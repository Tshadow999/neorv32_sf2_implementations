-- ********************************************************************/
-- Actel Corporation Proprietary and Confidential
--  Copyright 2011 Actel Corporation.  All rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
-- ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
-- IN ADVANCE IN WRITING.
--
-- Description:  SRAM block, 1 byte wide, 2048 to 141312 deep 
--              (in steps of 2048), used to construct the memory.
--
-- Revision Information:
-- Date     Description
--
-- SVN Revision Information:
-- SVN $Revision: 4805 $
-- SVN $Date: 2008-11-27 17:48:48 +0530 (Thu, 27 Nov 2008) $
--
-- Resolved SARs
-- SAR      Date     Who   Description
--
-- Notes:
--
-- ********************************************************************/
library ieee;
use     ieee.std_logic_1164.all;
use     ieee.std_logic_arith.all;
use     ieee.std_logic_unsigned.all;
use     ieee.std_logic_misc.all;
--use     work.XHDL_std_logic.all;
--use     work.XHDL_misc.all;


ENTITY COREAPBLSRAM_C0_COREAPBLSRAM_C0_0_lsram_2048to141312x8 IS
   GENERIC (
      -- ---------------------------------------------------------------------
      -- Parameters
      -- ---------------------------------------------------------------------
      -- DEPTH can range from 2048 to 141312, in steps of 2048
      DEPTH                          :  integer := 2048;    
      APB_DWIDTH                     :  integer := 8);    
   PORT (
      -- ---------------------------------------------------------------------
-- Port declarations
-- ---------------------------------------------------------------------
-- AhbFabric interface
-- Inputs

      writeData               : IN std_logic_vector(APB_DWIDTH - 1 
      DOWNTO 0);   
      -- Output

      readData                : OUT std_logic_vector(APB_DWIDTH - 1 
      DOWNTO 0);   
      -- AhbSramIf interface
-- Inputs

      wen                     : IN std_logic;   
      ren                     : IN std_logic;   
      writeAddr               : IN std_logic_vector(17 DOWNTO 0);   
      readAddr                : IN std_logic_vector(17 DOWNTO 0);   
      clk                     : IN std_logic;   
      resetn                  : IN std_logic;   
      lsram_2k_BUSY_all       : OUT std_logic);   
END ENTITY COREAPBLSRAM_C0_COREAPBLSRAM_C0_0_lsram_2048to141312x8;

ARCHITECTURE translated OF COREAPBLSRAM_C0_COREAPBLSRAM_C0_0_lsram_2048to141312x8 IS
   COMPONENT RAM1K18 
      PORT (
         A_DOUT               : OUT std_logic_vector(17 DOWNTO 0); 
         B_DOUT               : OUT std_logic_vector(17 DOWNTO 0); 
         A_CLK                : IN std_logic;
         B_CLK                : IN std_logic; 
         A_ARST_N                : IN std_logic; 
         B_ARST_N                 : IN std_logic;
         A_BLK              : IN std_logic_vector(2 DOWNTO 0);
         B_BLK              : IN std_logic_vector(2 DOWNTO 0);
         A_DIN              : IN std_logic_vector(17 DOWNTO 0);
         B_DIN              : IN std_logic_vector(17 DOWNTO 0);
         A_ADDR              : IN std_logic_vector(13 DOWNTO 0);
         B_ADDR              : IN std_logic_vector(13 DOWNTO 0);
         A_WEN              : IN std_logic_vector(1 DOWNTO 0);
         B_WEN              : IN std_logic_vector(1 DOWNTO 0);
         A_DOUT_CLK                : IN std_logic;
         B_DOUT_CLK                : IN std_logic;
         A_DOUT_EN                : IN std_logic;
         B_DOUT_EN                : IN std_logic;
         A_DOUT_ARST_N                : IN std_logic;
         B_DOUT_ARST_N                : IN std_logic;
         A_DOUT_SRST_N                : IN std_logic;
         B_DOUT_SRST_N                : IN std_logic;
         A_DOUT_LAT                : IN std_logic;
         B_DOUT_LAT                : IN std_logic;
         A_WIDTH              : IN std_logic_vector(2 DOWNTO 0);
         B_WIDTH              : IN std_logic_vector(2 DOWNTO 0);
         A_WMODE                : IN std_logic;
         B_WMODE                : IN std_logic;
         A_EN                : IN std_logic;
         B_EN                : IN std_logic;
         BUSY                : OUT std_logic;
         SII_LOCK                : IN std_logic);
  END COMPONENT;    


   -- ---------------------------------------------------------------------
   -- Constant declarations
   -- ---------------------------------------------------------------------
   -- ---------------------------------------------------------------------
   -- Signal declarations
   -- ---------------------------------------------------------------------
   SIGNAL ckRdAddr                 :  std_logic_vector(17 DOWNTO 9);   
   SIGNAL width0                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width1                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width2                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width3                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width4                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width5                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width6                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width7                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width8                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width9                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width10                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width11                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width12                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width13                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width14                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width15                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width16                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width17                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width18                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width19                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width20                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width21                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width22                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width23                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width24                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width25                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width26                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width27                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width28                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width29                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width30                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width31                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width32                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width33                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width34                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width35                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width36                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width37                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width38                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width39                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width40                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width41                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width42                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width43                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width44                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width45                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width46                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width47                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width48                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width49                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width50                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width51                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width52                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width53                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width54                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width55                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width56                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width57                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width58                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width59                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width60                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width61                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width62                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width63                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width64                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width65                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width66                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width67                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width68                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL wen_a0                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a1                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a2                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a3                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a4                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a5                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a6                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a7                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a8                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a9                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a10                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a11                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a12                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a13                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a14                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a15                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a16                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a17                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a18                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a19                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a20                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a21                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a22                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a23                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a24                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a25                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a26                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a27                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a28                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a29                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a30                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a31                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a32                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a33                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a34                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a35                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a36                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a37                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a38                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a39                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a40                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a41                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a42                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a43                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a44                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a45                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a46                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a47                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a48                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a49                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a50                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a51                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a52                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a53                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a54                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a55                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a56                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a57                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a58                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a59                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a60                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a61                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a62                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a63                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a64                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a65                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a66                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a67                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_a68                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b0                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b1                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b2                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b3                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b4                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b5                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b6                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b7                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b8                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b9                   :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b10                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b11                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b12                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b13                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b14                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b15                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b16                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b17                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b18                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b19                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b20                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b21                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b22                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b23                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b24                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b25                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b26                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b27                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b28                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b29                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b30                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b31                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b32                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b33                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b34                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b35                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b36                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b37                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b38                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b39                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b40                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b41                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b42                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b43                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b44                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b45                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b46                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b47                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b48                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b49                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b50                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b51                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b52                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b53                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b54                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b55                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b56                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b57                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b58                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b59                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b60                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b61                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b62                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b63                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b64                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b65                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b66                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b67                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL wen_b68                  :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL writeData0               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData1               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData2               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData3               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData4               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData5               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData6               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData7               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData8               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData9               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData10              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData11              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData12              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData13              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData14              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData15              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData16              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData17              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData18              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData19              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData20              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData21              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData22              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData23              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData24              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData25              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData26              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData27              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData28              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData29              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData30              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData31              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData32              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData33              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData34              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData35              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData36              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData37              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData38              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData39              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData40              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData41              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData42              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData43              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData44              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData45              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData46              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData47              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData48              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData49              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData50              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData51              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData52              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData53              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData54              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData55              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData56              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData57              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData58              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData59              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData60              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData61              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData62              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData63              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData64              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData65              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData66              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData67              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData68              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData0                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData1                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData2                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData3                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData4                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData5                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData6                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData7                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData8                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData9                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData10               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData11               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData12               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData13               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData14               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData15               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData16               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData17               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData18               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData19               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData20               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData21               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData22               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData23               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData24               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData25               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData26               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData27               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData28               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData29               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData30               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData31               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData32               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData33               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData34               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData35               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData36               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData37               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData38               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData39               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData40               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData41               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData42               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData43               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData44               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData45               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData46               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData47               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData48               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData49               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData50               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData51               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData52               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData53               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData54               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData55               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData56               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData57               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData58               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData59               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData60               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData61               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData62               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData63               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData64               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData65               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData66               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData67               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData68               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeAddr0               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr1               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr2               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr3               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr4               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr5               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr6               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr7               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr8               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr9               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr10              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr11              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr12              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr13              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr14              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr15              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr16              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr17              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr18              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr19              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr20              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr21              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr22              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr23              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr24              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr25              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr26              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr27              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr28              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr29              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr30              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr31              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr32              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr33              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr34              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr35              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr36              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr37              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr38              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr39              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr40              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr41              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr42              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr43              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr44              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr45              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr46              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr47              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr48              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr49              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr50              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr51              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr52              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr53              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr54              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr55              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr56              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr57              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr58              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr59              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr60              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr61              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr62              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr63              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr64              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr65              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr66              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr67              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL writeAddr68              :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr0                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr1                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr2                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr3                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr4                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr5                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr6                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr7                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr8                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr9                :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr10               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr11               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr12               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr13               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr14               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr15               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr16               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr17               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr18               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr19               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr20               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr21               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr22               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr23               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr24               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr25               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr26               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr27               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr28               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr29               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr30               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr31               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr32               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr33               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr34               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr35               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr36               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr37               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr38               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr39               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr40               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr41               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr42               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr43               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr44               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr45               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr46               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr47               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr48               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr49               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr50               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr51               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr52               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr53               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr54               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr55               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr56               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr57               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr58               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr59               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr60               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr61               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr62               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr63               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr64               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr65               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr66               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr67               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL readAddr68               :  std_logic_vector(13 DOWNTO 0);   
   SIGNAL lsram_2k_BUSY_68         :  std_logic;   
   SIGNAL lsram_2k_BUSY_67         :  std_logic;   
   SIGNAL lsram_2k_BUSY_66         :  std_logic;   
   SIGNAL lsram_2k_BUSY_65         :  std_logic;   
   SIGNAL lsram_2k_BUSY_64         :  std_logic;   
   SIGNAL lsram_2k_BUSY_63         :  std_logic;   
   SIGNAL lsram_2k_BUSY_62         :  std_logic;   
   SIGNAL lsram_2k_BUSY_61         :  std_logic;   
   SIGNAL lsram_2k_BUSY_60         :  std_logic;   
   SIGNAL lsram_2k_BUSY_59         :  std_logic;   
   SIGNAL lsram_2k_BUSY_58         :  std_logic;   
   SIGNAL lsram_2k_BUSY_57         :  std_logic;   
   SIGNAL lsram_2k_BUSY_56         :  std_logic;   
   SIGNAL lsram_2k_BUSY_55         :  std_logic;   
   SIGNAL lsram_2k_BUSY_54         :  std_logic;   
   SIGNAL lsram_2k_BUSY_53         :  std_logic;   
   SIGNAL lsram_2k_BUSY_52         :  std_logic;   
   SIGNAL lsram_2k_BUSY_51         :  std_logic;   
   SIGNAL lsram_2k_BUSY_50         :  std_logic;   
   SIGNAL lsram_2k_BUSY_49         :  std_logic;   
   SIGNAL lsram_2k_BUSY_48         :  std_logic;   
   SIGNAL lsram_2k_BUSY_47         :  std_logic;   
   SIGNAL lsram_2k_BUSY_46         :  std_logic;   
   SIGNAL lsram_2k_BUSY_45         :  std_logic;   
   SIGNAL lsram_2k_BUSY_44         :  std_logic;   
   SIGNAL lsram_2k_BUSY_43         :  std_logic;   
   SIGNAL lsram_2k_BUSY_42         :  std_logic;   
   SIGNAL lsram_2k_BUSY_41         :  std_logic;   
   SIGNAL lsram_2k_BUSY_40         :  std_logic;   
   SIGNAL lsram_2k_BUSY_39         :  std_logic;   
   SIGNAL lsram_2k_BUSY_38         :  std_logic;   
   SIGNAL lsram_2k_BUSY_37         :  std_logic;   
   SIGNAL lsram_2k_BUSY_36         :  std_logic;   
   SIGNAL lsram_2k_BUSY_35         :  std_logic;   
   SIGNAL lsram_2k_BUSY_34         :  std_logic;   
   SIGNAL lsram_2k_BUSY_33         :  std_logic;   
   SIGNAL lsram_2k_BUSY_32         :  std_logic;   
   SIGNAL lsram_2k_BUSY_31         :  std_logic;   
   SIGNAL lsram_2k_BUSY_30         :  std_logic;   
   SIGNAL lsram_2k_BUSY_29         :  std_logic;   
   SIGNAL lsram_2k_BUSY_28         :  std_logic;   
   SIGNAL lsram_2k_BUSY_27         :  std_logic;   
   SIGNAL lsram_2k_BUSY_26         :  std_logic;   
   SIGNAL lsram_2k_BUSY_25         :  std_logic;   
   SIGNAL lsram_2k_BUSY_24         :  std_logic;   
   SIGNAL lsram_2k_BUSY_23         :  std_logic;   
   SIGNAL lsram_2k_BUSY_22         :  std_logic;   
   SIGNAL lsram_2k_BUSY_21         :  std_logic;   
   SIGNAL lsram_2k_BUSY_20         :  std_logic;   
   SIGNAL lsram_2k_BUSY_19         :  std_logic;   
   SIGNAL lsram_2k_BUSY_18         :  std_logic;   
   SIGNAL lsram_2k_BUSY_17         :  std_logic;   
   SIGNAL lsram_2k_BUSY_16         :  std_logic;   
   SIGNAL lsram_2k_BUSY_15         :  std_logic;   
   SIGNAL lsram_2k_BUSY_14         :  std_logic;   
   SIGNAL lsram_2k_BUSY_13         :  std_logic;   
   SIGNAL lsram_2k_BUSY_12         :  std_logic;   
   SIGNAL lsram_2k_BUSY_11         :  std_logic;   
   SIGNAL lsram_2k_BUSY_10         :  std_logic;   
   SIGNAL lsram_2k_BUSY_9          :  std_logic;   
   SIGNAL lsram_2k_BUSY_8          :  std_logic;   
   SIGNAL lsram_2k_BUSY_7          :  std_logic;   
   SIGNAL lsram_2k_BUSY_6          :  std_logic;   
   SIGNAL lsram_2k_BUSY_5          :  std_logic;   
   SIGNAL lsram_2k_BUSY_4          :  std_logic;   
   SIGNAL lsram_2k_BUSY_3          :  std_logic;   
   SIGNAL lsram_2k_BUSY_2          :  std_logic;   
   SIGNAL lsram_2k_BUSY_1          :  std_logic;   
   SIGNAL lsram_2k_BUSY_0          :  std_logic;   
   SIGNAL readData_xhdl1           :  std_logic_vector(APB_DWIDTH - 1 
   DOWNTO 0);   
   SIGNAL lsram_2k_BUSY_all_xhdl2  :  std_logic;   

BEGIN
   readData <= readData_xhdl1;
   lsram_2k_BUSY_all <= lsram_2k_BUSY_all_xhdl2;

   ------------------------------------------------------------------------
   -- Main body of code
   ------------------------------------------------------------------------
   
   PROCESS (clk, resetn)
   BEGIN
      IF (NOT resetn = '1') THEN
         ckRdAddr(17 DOWNTO 9) <= "000000000";    
      ELSIF (clk'EVENT AND clk = '1') THEN
         ckRdAddr(17 DOWNTO 9) <= readAddr(17 DOWNTO 9);    
      END IF;
   END PROCESS;

   ------------------------------------------------------------------------------------------
   -- Assign values to various signals based on DEPTH and RAM4K9_WIDTH settings.
   -- Default is to build the (byte wide) memory from RAM blocks which are configured to
   -- be tall and narrow.
   ------------------------------------------------------------------------------------------
   
   PROCESS (readData20, readData21, readData22, readData23, readData24, 
   readData25, readData26, readData27, readData60, readData61, 
   readData28, readData62, readData29, readData63, readData64, 
   readData65, readData66, readData67, readData68, clk, 
   readData30, readData31, writeData, readData32, readData33, resetn, 
   readData34, readData35, readData36, readData37, readData38, 
   readData39, ckRdAddr, readData40, readData41, readData42, 
   readData43, readData44, readData45, readAddr, readData46, readData47, 
   readData48, readData49, readData10, readData11, readData12, 
   readData13, readData14, readData15, wen, readData16, readData17, 
   readData0, readData50, readData18, readData1, readData51, readData2, 
   readData52, readData19, readData3, readData53, readData4, readData54, 
   readData5, readData6, readData55, readData7, readData56, readData8, 
   readData57, readData9, readData58, readData59, writeAddr)
      VARIABLE width0_xhdl3  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width1_xhdl4  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width2_xhdl5  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width3_xhdl6  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width4_xhdl7  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width5_xhdl8  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width6_xhdl9  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width7_xhdl10  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width8_xhdl11  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width9_xhdl12  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width10_xhdl13  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width11_xhdl14  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width12_xhdl15  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width13_xhdl16  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width14_xhdl17  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width15_xhdl18  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width16_xhdl19  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width17_xhdl20  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width18_xhdl21  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width19_xhdl22  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width20_xhdl23  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width21_xhdl24  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width22_xhdl25  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width23_xhdl26  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width24_xhdl27  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width25_xhdl28  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width26_xhdl29  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width27_xhdl30  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width28_xhdl31  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width29_xhdl32  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width30_xhdl33  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width31_xhdl34  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width32_xhdl35  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width33_xhdl36  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width34_xhdl37  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width35_xhdl38  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width36_xhdl39  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width37_xhdl40  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width38_xhdl41  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width39_xhdl42  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width40_xhdl43  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width41_xhdl44  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width42_xhdl45  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width43_xhdl46  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width44_xhdl47  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width45_xhdl48  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width46_xhdl49  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width47_xhdl50  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width48_xhdl51  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width49_xhdl52  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width50_xhdl53  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width51_xhdl54  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width52_xhdl55  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width53_xhdl56  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width54_xhdl57  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width55_xhdl58  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width56_xhdl59  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width57_xhdl60  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width58_xhdl61  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width59_xhdl62  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width60_xhdl63  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width61_xhdl64  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width62_xhdl65  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width63_xhdl66  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width64_xhdl67  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width65_xhdl68  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width66_xhdl69  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width67_xhdl70  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width68_xhdl71  : std_logic_vector(2 DOWNTO 0);
      VARIABLE wen_a0_xhdl72  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a1_xhdl73  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a2_xhdl74  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a3_xhdl75  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a4_xhdl76  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a5_xhdl77  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a6_xhdl78  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a7_xhdl79  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a8_xhdl80  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a9_xhdl81  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a10_xhdl82  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a11_xhdl83  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a12_xhdl84  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a13_xhdl85  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a14_xhdl86  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a15_xhdl87  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a16_xhdl88  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a17_xhdl89  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a18_xhdl90  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a19_xhdl91  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a20_xhdl92  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a21_xhdl93  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a22_xhdl94  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a23_xhdl95  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a24_xhdl96  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a25_xhdl97  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a26_xhdl98  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a27_xhdl99  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a28_xhdl100  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a29_xhdl101  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a30_xhdl102  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a31_xhdl103  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a32_xhdl104  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a33_xhdl105  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a34_xhdl106  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a35_xhdl107  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a36_xhdl108  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a37_xhdl109  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a38_xhdl110  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a39_xhdl111  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a40_xhdl112  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a41_xhdl113  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a42_xhdl114  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a43_xhdl115  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a44_xhdl116  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a45_xhdl117  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a46_xhdl118  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a47_xhdl119  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a48_xhdl120  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a49_xhdl121  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a50_xhdl122  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a51_xhdl123  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a52_xhdl124  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a53_xhdl125  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a54_xhdl126  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a55_xhdl127  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a56_xhdl128  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a57_xhdl129  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a58_xhdl130  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a59_xhdl131  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a60_xhdl132  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a61_xhdl133  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a62_xhdl134  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a63_xhdl135  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a64_xhdl136  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a65_xhdl137  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a66_xhdl138  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a67_xhdl139  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_a68_xhdl140  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b0_xhdl141  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b1_xhdl142  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b2_xhdl143  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b3_xhdl144  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b4_xhdl145  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b5_xhdl146  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b6_xhdl147  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b7_xhdl148  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b8_xhdl149  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b9_xhdl150  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b10_xhdl151  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b11_xhdl152  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b12_xhdl153  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b13_xhdl154  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b14_xhdl155  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b15_xhdl156  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b16_xhdl157  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b17_xhdl158  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b18_xhdl159  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b19_xhdl160  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b20_xhdl161  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b21_xhdl162  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b22_xhdl163  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b23_xhdl164  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b24_xhdl165  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b25_xhdl166  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b26_xhdl167  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b27_xhdl168  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b28_xhdl169  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b29_xhdl170  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b30_xhdl171  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b31_xhdl172  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b32_xhdl173  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b33_xhdl174  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b34_xhdl175  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b35_xhdl176  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b36_xhdl177  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b37_xhdl178  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b38_xhdl179  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b39_xhdl180  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b40_xhdl181  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b41_xhdl182  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b42_xhdl183  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b43_xhdl184  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b44_xhdl185  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b45_xhdl186  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b46_xhdl187  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b47_xhdl188  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b48_xhdl189  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b49_xhdl190  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b50_xhdl191  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b51_xhdl192  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b52_xhdl193  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b53_xhdl194  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b54_xhdl195  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b55_xhdl196  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b56_xhdl197  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b57_xhdl198  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b58_xhdl199  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b59_xhdl200  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b60_xhdl201  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b61_xhdl202  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b62_xhdl203  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b63_xhdl204  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b64_xhdl205  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b65_xhdl206  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b66_xhdl207  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b67_xhdl208  : std_logic_vector(1 DOWNTO 0);
      VARIABLE wen_b68_xhdl209  : std_logic_vector(1 DOWNTO 0);
      VARIABLE writeData0_xhdl210  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData1_xhdl211  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData2_xhdl212  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData3_xhdl213  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData4_xhdl214  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData5_xhdl215  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData6_xhdl216  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData7_xhdl217  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData8_xhdl218  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData9_xhdl219  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData10_xhdl220  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData11_xhdl221  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData12_xhdl222  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData13_xhdl223  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData14_xhdl224  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData15_xhdl225  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData16_xhdl226  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData17_xhdl227  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData18_xhdl228  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData19_xhdl229  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData20_xhdl230  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData21_xhdl231  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData22_xhdl232  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData23_xhdl233  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData24_xhdl234  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData25_xhdl235  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData26_xhdl236  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData27_xhdl237  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData28_xhdl238  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData29_xhdl239  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData30_xhdl240  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData31_xhdl241  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData32_xhdl242  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData33_xhdl243  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData34_xhdl244  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData35_xhdl245  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData36_xhdl246  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData37_xhdl247  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData38_xhdl248  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData39_xhdl249  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData40_xhdl250  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData41_xhdl251  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData42_xhdl252  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData43_xhdl253  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData44_xhdl254  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData45_xhdl255  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData46_xhdl256  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData47_xhdl257  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData48_xhdl258  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData49_xhdl259  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData50_xhdl260  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData51_xhdl261  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData52_xhdl262  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData53_xhdl263  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData54_xhdl264  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData55_xhdl265  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData56_xhdl266  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData57_xhdl267  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData58_xhdl268  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData59_xhdl269  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData60_xhdl270  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData61_xhdl271  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData62_xhdl272  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData63_xhdl273  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData64_xhdl274  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData65_xhdl275  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData66_xhdl276  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData67_xhdl277  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData68_xhdl278  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeAddr0_xhdl279  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr1_xhdl280  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr2_xhdl281  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr3_xhdl282  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr4_xhdl283  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr5_xhdl284  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr6_xhdl285  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr7_xhdl286  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr8_xhdl287  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr9_xhdl288  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr10_xhdl289  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr11_xhdl290  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr12_xhdl291  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr13_xhdl292  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr14_xhdl293  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr15_xhdl294  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr16_xhdl295  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr17_xhdl296  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr18_xhdl297  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr19_xhdl298  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr20_xhdl299  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr21_xhdl300  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr22_xhdl301  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr23_xhdl302  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr24_xhdl303  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr25_xhdl304  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr26_xhdl305  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr27_xhdl306  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr28_xhdl307  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr29_xhdl308  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr30_xhdl309  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr31_xhdl310  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr32_xhdl311  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr33_xhdl312  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr34_xhdl313  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr35_xhdl314  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr36_xhdl315  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr37_xhdl316  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr38_xhdl317  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr39_xhdl318  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr40_xhdl319  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr41_xhdl320  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr42_xhdl321  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr43_xhdl322  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr44_xhdl323  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr45_xhdl324  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr46_xhdl325  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr47_xhdl326  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr48_xhdl327  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr49_xhdl328  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr50_xhdl329  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr51_xhdl330  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr52_xhdl331  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr53_xhdl332  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr54_xhdl333  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr55_xhdl334  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr56_xhdl335  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr57_xhdl336  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr58_xhdl337  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr59_xhdl338  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr60_xhdl339  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr61_xhdl340  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr62_xhdl341  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr63_xhdl342  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr64_xhdl343  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr65_xhdl344  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr66_xhdl345  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr67_xhdl346  : std_logic_vector(13 DOWNTO 0);
      VARIABLE writeAddr68_xhdl347  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr0_xhdl348  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr1_xhdl349  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr2_xhdl350  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr3_xhdl351  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr4_xhdl352  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr5_xhdl353  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr6_xhdl354  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr7_xhdl355  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr8_xhdl356  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr9_xhdl357  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr10_xhdl358  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr11_xhdl359  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr12_xhdl360  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr13_xhdl361  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr14_xhdl362  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr15_xhdl363  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr16_xhdl364  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr17_xhdl365  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr18_xhdl366  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr19_xhdl367  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr20_xhdl368  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr21_xhdl369  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr22_xhdl370  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr23_xhdl371  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr24_xhdl372  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr25_xhdl373  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr26_xhdl374  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr27_xhdl375  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr28_xhdl376  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr29_xhdl377  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr30_xhdl378  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr31_xhdl379  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr32_xhdl380  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr33_xhdl381  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr34_xhdl382  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr35_xhdl383  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr36_xhdl384  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr37_xhdl385  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr38_xhdl386  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr39_xhdl387  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr40_xhdl388  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr41_xhdl389  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr42_xhdl390  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr43_xhdl391  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr44_xhdl392  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr45_xhdl393  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr46_xhdl394  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr47_xhdl395  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr48_xhdl396  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr49_xhdl397  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr50_xhdl398  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr51_xhdl399  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr52_xhdl400  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr53_xhdl401  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr54_xhdl402  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr55_xhdl403  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr56_xhdl404  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr57_xhdl405  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr58_xhdl406  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr59_xhdl407  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr60_xhdl408  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr61_xhdl409  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr62_xhdl410  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr63_xhdl411  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr64_xhdl412  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr65_xhdl413  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr66_xhdl414  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr67_xhdl415  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readAddr68_xhdl416  : std_logic_vector(13 DOWNTO 0);
      VARIABLE readData_xhdl1_xhdl417  : std_logic_vector(APB_DWIDTH - 1 
      DOWNTO 0);
   BEGIN
      width0_xhdl3 := "000";    
      width1_xhdl4 := "000";    
      width2_xhdl5 := "000";    
      width3_xhdl6 := "000";    
      width4_xhdl7 := "000";    
      width5_xhdl8 := "000";    
      width6_xhdl9 := "000";    
      width7_xhdl10 := "000";    
      width8_xhdl11 := "000";    
      width9_xhdl12 := "000";    
      width10_xhdl13 := "000";    
      width11_xhdl14 := "000";    
      width12_xhdl15 := "000";    
      width13_xhdl16 := "000";    
      width14_xhdl17 := "000";    
      width15_xhdl18 := "000";    
      width16_xhdl19 := "000";    
      width17_xhdl20 := "000";    
      width18_xhdl21 := "000";    
      width19_xhdl22 := "000";    
      width20_xhdl23 := "000";    
      width21_xhdl24 := "000";    
      width22_xhdl25 := "000";    
      width23_xhdl26 := "000";    
      width24_xhdl27 := "000";    
      width25_xhdl28 := "000";    
      width26_xhdl29 := "000";    
      width27_xhdl30 := "000";    
      width28_xhdl31 := "000";    
      width29_xhdl32 := "000";    
      width30_xhdl33 := "000";    
      width31_xhdl34 := "000";    
      width32_xhdl35 := "000";    
      width33_xhdl36 := "000";    
      width34_xhdl37 := "000";    
      width35_xhdl38 := "000";    
      width36_xhdl39 := "000";    
      width37_xhdl40 := "000";    
      width38_xhdl41 := "000";    
      width39_xhdl42 := "000";    
      width40_xhdl43 := "000";    
      width41_xhdl44 := "000";    
      width42_xhdl45 := "000";    
      width43_xhdl46 := "000";    
      width44_xhdl47 := "000";    
      width45_xhdl48 := "000";    
      width46_xhdl49 := "000";    
      width47_xhdl50 := "000";    
      width48_xhdl51 := "000";    
      width49_xhdl52 := "000";    
      width50_xhdl53 := "000";    
      width51_xhdl54 := "000";    
      width52_xhdl55 := "000";    
      width53_xhdl56 := "000";    
      width54_xhdl57 := "000";    
      width55_xhdl58 := "000";    
      width56_xhdl59 := "000";    
      width57_xhdl60 := "000";    
      width58_xhdl61 := "000";    
      width59_xhdl62 := "000";    
      width60_xhdl63 := "000";    
      width61_xhdl64 := "000";    
      width62_xhdl65 := "000";    
      width63_xhdl66 := "000";    
      width64_xhdl67 := "000";    
      width65_xhdl68 := "000";    
      width66_xhdl69 := "000";    
      width67_xhdl70 := "000";    
      width68_xhdl71 := "000";    
      wen_a0_xhdl72 := "00";    
      wen_a1_xhdl73 := "00";    
      wen_a2_xhdl74 := "00";    
      wen_a3_xhdl75 := "00";    
      wen_a4_xhdl76 := "00";    
      wen_a5_xhdl77 := "00";    
      wen_a6_xhdl78 := "00";    
      wen_a7_xhdl79 := "00";    
      wen_a8_xhdl80 := "00";    
      wen_a9_xhdl81 := "00";    
      wen_a10_xhdl82 := "00";    
      wen_a11_xhdl83 := "00";    
      wen_a12_xhdl84 := "00";    
      wen_a13_xhdl85 := "00";    
      wen_a14_xhdl86 := "00";    
      wen_a15_xhdl87 := "00";    
      wen_a16_xhdl88 := "00";    
      wen_a17_xhdl89 := "00";    
      wen_a18_xhdl90 := "00";    
      wen_a19_xhdl91 := "00";    
      wen_a20_xhdl92 := "00";    
      wen_a21_xhdl93 := "00";    
      wen_a22_xhdl94 := "00";    
      wen_a23_xhdl95 := "00";    
      wen_a24_xhdl96 := "00";    
      wen_a25_xhdl97 := "00";    
      wen_a26_xhdl98 := "00";    
      wen_a27_xhdl99 := "00";    
      wen_a28_xhdl100 := "00";    
      wen_a29_xhdl101 := "00";    
      wen_a30_xhdl102 := "00";    
      wen_a31_xhdl103 := "00";    
      wen_a32_xhdl104 := "00";    
      wen_a33_xhdl105 := "00";    
      wen_a34_xhdl106 := "00";    
      wen_a35_xhdl107 := "00";    
      wen_a36_xhdl108 := "00";    
      wen_a37_xhdl109 := "00";    
      wen_a38_xhdl110 := "00";    
      wen_a39_xhdl111 := "00";    
      wen_a40_xhdl112 := "00";    
      wen_a41_xhdl113 := "00";    
      wen_a42_xhdl114 := "00";    
      wen_a43_xhdl115 := "00";    
      wen_a44_xhdl116 := "00";    
      wen_a45_xhdl117 := "00";    
      wen_a46_xhdl118 := "00";    
      wen_a47_xhdl119 := "00";    
      wen_a48_xhdl120 := "00";    
      wen_a49_xhdl121 := "00";    
      wen_a50_xhdl122 := "00";    
      wen_a51_xhdl123 := "00";    
      wen_a52_xhdl124 := "00";    
      wen_a53_xhdl125 := "00";    
      wen_a54_xhdl126 := "00";    
      wen_a55_xhdl127 := "00";    
      wen_a56_xhdl128 := "00";    
      wen_a57_xhdl129 := "00";    
      wen_a58_xhdl130 := "00";    
      wen_a59_xhdl131 := "00";    
      wen_a60_xhdl132 := "00";    
      wen_a61_xhdl133 := "00";    
      wen_a62_xhdl134 := "00";    
      wen_a63_xhdl135 := "00";    
      wen_a64_xhdl136 := "00";    
      wen_a65_xhdl137 := "00";    
      wen_a66_xhdl138 := "00";    
      wen_a67_xhdl139 := "00";    
      wen_a68_xhdl140 := "00";    
      wen_b0_xhdl141 := "00";    
      wen_b1_xhdl142 := "00";    
      wen_b2_xhdl143 := "00";    
      wen_b3_xhdl144 := "00";    
      wen_b4_xhdl145 := "00";    
      wen_b5_xhdl146 := "00";    
      wen_b6_xhdl147 := "00";    
      wen_b7_xhdl148 := "00";    
      wen_b8_xhdl149 := "00";    
      wen_b9_xhdl150 := "00";    
      wen_b10_xhdl151 := "00";    
      wen_b11_xhdl152 := "00";    
      wen_b12_xhdl153 := "00";    
      wen_b13_xhdl154 := "00";    
      wen_b14_xhdl155 := "00";    
      wen_b15_xhdl156 := "00";    
      wen_b16_xhdl157 := "00";    
      wen_b17_xhdl158 := "00";    
      wen_b18_xhdl159 := "00";    
      wen_b19_xhdl160 := "00";    
      wen_b20_xhdl161 := "00";    
      wen_b21_xhdl162 := "00";    
      wen_b22_xhdl163 := "00";    
      wen_b23_xhdl164 := "00";    
      wen_b24_xhdl165 := "00";    
      wen_b25_xhdl166 := "00";    
      wen_b26_xhdl167 := "00";    
      wen_b27_xhdl168 := "00";    
      wen_b28_xhdl169 := "00";    
      wen_b29_xhdl170 := "00";    
      wen_b30_xhdl171 := "00";    
      wen_b31_xhdl172 := "00";    
      wen_b32_xhdl173 := "00";    
      wen_b33_xhdl174 := "00";    
      wen_b34_xhdl175 := "00";    
      wen_b35_xhdl176 := "00";    
      wen_b36_xhdl177 := "00";    
      wen_b37_xhdl178 := "00";    
      wen_b38_xhdl179 := "00";    
      wen_b39_xhdl180 := "00";    
      wen_b40_xhdl181 := "00";    
      wen_b41_xhdl182 := "00";    
      wen_b42_xhdl183 := "00";    
      wen_b43_xhdl184 := "00";    
      wen_b44_xhdl185 := "00";    
      wen_b45_xhdl186 := "00";    
      wen_b46_xhdl187 := "00";    
      wen_b47_xhdl188 := "00";    
      wen_b48_xhdl189 := "00";    
      wen_b49_xhdl190 := "00";    
      wen_b50_xhdl191 := "00";    
      wen_b51_xhdl192 := "00";    
      wen_b52_xhdl193 := "00";    
      wen_b53_xhdl194 := "00";    
      wen_b54_xhdl195 := "00";    
      wen_b55_xhdl196 := "00";    
      wen_b56_xhdl197 := "00";    
      wen_b57_xhdl198 := "00";    
      wen_b58_xhdl199 := "00";    
      wen_b59_xhdl200 := "00";    
      wen_b60_xhdl201 := "00";    
      wen_b61_xhdl202 := "00";    
      wen_b62_xhdl203 := "00";    
      wen_b63_xhdl204 := "00";    
      wen_b64_xhdl205 := "00";    
      wen_b65_xhdl206 := "00";    
      wen_b66_xhdl207 := "00";    
      wen_b67_xhdl208 := "00";    
      wen_b68_xhdl209 := "00";    
      writeData0_xhdl210 := "000000000000000000";    
      writeData1_xhdl211 := "000000000000000000";    
      writeData2_xhdl212 := "000000000000000000";    
      writeData3_xhdl213 := "000000000000000000";    
      writeData4_xhdl214 := "000000000000000000";    
      writeData5_xhdl215 := "000000000000000000";    
      writeData6_xhdl216 := "000000000000000000";    
      writeData7_xhdl217 := "000000000000000000";    
      writeData8_xhdl218 := "000000000000000000";    
      writeData9_xhdl219 := "000000000000000000";    
      writeData10_xhdl220 := "000000000000000000";    
      writeData11_xhdl221 := "000000000000000000";    
      writeData12_xhdl222 := "000000000000000000";    
      writeData13_xhdl223 := "000000000000000000";    
      writeData14_xhdl224 := "000000000000000000";    
      writeData15_xhdl225 := "000000000000000000";    
      writeData16_xhdl226 := "000000000000000000";    
      writeData17_xhdl227 := "000000000000000000";    
      writeData18_xhdl228 := "000000000000000000";    
      writeData19_xhdl229 := "000000000000000000";    
      writeData20_xhdl230 := "000000000000000000";    
      writeData21_xhdl231 := "000000000000000000";    
      writeData22_xhdl232 := "000000000000000000";    
      writeData23_xhdl233 := "000000000000000000";    
      writeData24_xhdl234 := "000000000000000000";    
      writeData25_xhdl235 := "000000000000000000";    
      writeData26_xhdl236 := "000000000000000000";    
      writeData27_xhdl237 := "000000000000000000";    
      writeData28_xhdl238 := "000000000000000000";    
      writeData29_xhdl239 := "000000000000000000";    
      writeData30_xhdl240 := "000000000000000000";    
      writeData31_xhdl241 := "000000000000000000";    
      writeData32_xhdl242 := "000000000000000000";    
      writeData33_xhdl243 := "000000000000000000";    
      writeData34_xhdl244 := "000000000000000000";    
      writeData35_xhdl245 := "000000000000000000";    
      writeData36_xhdl246 := "000000000000000000";    
      writeData37_xhdl247 := "000000000000000000";    
      writeData38_xhdl248 := "000000000000000000";    
      writeData39_xhdl249 := "000000000000000000";    
      writeData40_xhdl250 := "000000000000000000";    
      writeData41_xhdl251 := "000000000000000000";    
      writeData42_xhdl252 := "000000000000000000";    
      writeData43_xhdl253 := "000000000000000000";    
      writeData44_xhdl254 := "000000000000000000";    
      writeData45_xhdl255 := "000000000000000000";    
      writeData46_xhdl256 := "000000000000000000";    
      writeData47_xhdl257 := "000000000000000000";    
      writeData48_xhdl258 := "000000000000000000";    
      writeData49_xhdl259 := "000000000000000000";    
      writeData50_xhdl260 := "000000000000000000";    
      writeData51_xhdl261 := "000000000000000000";    
      writeData52_xhdl262 := "000000000000000000";    
      writeData53_xhdl263 := "000000000000000000";    
      writeData54_xhdl264 := "000000000000000000";    
      writeData55_xhdl265 := "000000000000000000";    
      writeData56_xhdl266 := "000000000000000000";    
      writeData57_xhdl267 := "000000000000000000";    
      writeData58_xhdl268 := "000000000000000000";    
      writeData59_xhdl269 := "000000000000000000";    
      writeData60_xhdl270 := "000000000000000000";    
      writeData61_xhdl271 := "000000000000000000";    
      writeData62_xhdl272 := "000000000000000000";    
      writeData63_xhdl273 := "000000000000000000";    
      writeData64_xhdl274 := "000000000000000000";    
      writeData65_xhdl275 := "000000000000000000";    
      writeData66_xhdl276 := "000000000000000000";    
      writeData67_xhdl277 := "000000000000000000";    
      writeData68_xhdl278 := "000000000000000000";    
      writeAddr0_xhdl279 := "00000000000000";    
      writeAddr1_xhdl280 := "00000000000000";    
      writeAddr2_xhdl281 := "00000000000000";    
      writeAddr3_xhdl282 := "00000000000000";    
      writeAddr4_xhdl283 := "00000000000000";    
      writeAddr5_xhdl284 := "00000000000000";    
      writeAddr6_xhdl285 := "00000000000000";    
      writeAddr7_xhdl286 := "00000000000000";    
      writeAddr8_xhdl287 := "00000000000000";    
      writeAddr9_xhdl288 := "00000000000000";    
      writeAddr10_xhdl289 := "00000000000000";    
      writeAddr11_xhdl290 := "00000000000000";    
      writeAddr12_xhdl291 := "00000000000000";    
      writeAddr13_xhdl292 := "00000000000000";    
      writeAddr14_xhdl293 := "00000000000000";    
      writeAddr15_xhdl294 := "00000000000000";    
      writeAddr16_xhdl295 := "00000000000000";    
      writeAddr17_xhdl296 := "00000000000000";    
      writeAddr18_xhdl297 := "00000000000000";    
      writeAddr19_xhdl298 := "00000000000000";    
      writeAddr20_xhdl299 := "00000000000000";    
      writeAddr21_xhdl300 := "00000000000000";    
      writeAddr22_xhdl301 := "00000000000000";    
      writeAddr23_xhdl302 := "00000000000000";    
      writeAddr24_xhdl303 := "00000000000000";    
      writeAddr25_xhdl304 := "00000000000000";    
      writeAddr26_xhdl305 := "00000000000000";    
      writeAddr27_xhdl306 := "00000000000000";    
      writeAddr28_xhdl307 := "00000000000000";    
      writeAddr29_xhdl308 := "00000000000000";    
      writeAddr30_xhdl309 := "00000000000000";    
      writeAddr31_xhdl310 := "00000000000000";    
      writeAddr32_xhdl311 := "00000000000000";    
      writeAddr33_xhdl312 := "00000000000000";    
      writeAddr34_xhdl313 := "00000000000000";    
      writeAddr35_xhdl314 := "00000000000000";    
      writeAddr36_xhdl315 := "00000000000000";    
      writeAddr37_xhdl316 := "00000000000000";    
      writeAddr38_xhdl317 := "00000000000000";    
      writeAddr39_xhdl318 := "00000000000000";    
      writeAddr40_xhdl319 := "00000000000000";    
      writeAddr41_xhdl320 := "00000000000000";    
      writeAddr42_xhdl321 := "00000000000000";    
      writeAddr43_xhdl322 := "00000000000000";    
      writeAddr44_xhdl323 := "00000000000000";    
      writeAddr45_xhdl324 := "00000000000000";    
      writeAddr46_xhdl325 := "00000000000000";    
      writeAddr47_xhdl326 := "00000000000000";    
      writeAddr48_xhdl327 := "00000000000000";    
      writeAddr49_xhdl328 := "00000000000000";    
      writeAddr50_xhdl329 := "00000000000000";    
      writeAddr51_xhdl330 := "00000000000000";    
      writeAddr52_xhdl331 := "00000000000000";    
      writeAddr53_xhdl332 := "00000000000000";    
      writeAddr54_xhdl333 := "00000000000000";    
      writeAddr55_xhdl334 := "00000000000000";    
      writeAddr56_xhdl335 := "00000000000000";    
      writeAddr57_xhdl336 := "00000000000000";    
      writeAddr58_xhdl337 := "00000000000000";    
      writeAddr59_xhdl338 := "00000000000000";    
      writeAddr60_xhdl339 := "00000000000000";    
      writeAddr61_xhdl340 := "00000000000000";    
      writeAddr62_xhdl341 := "00000000000000";    
      writeAddr63_xhdl342 := "00000000000000";    
      writeAddr64_xhdl343 := "00000000000000";    
      writeAddr65_xhdl344 := "00000000000000";    
      writeAddr66_xhdl345 := "00000000000000";    
      writeAddr67_xhdl346 := "00000000000000";    
      writeAddr68_xhdl347 := "00000000000000";    
      readAddr0_xhdl348 := "00000000000000";    
      readAddr1_xhdl349 := "00000000000000";    
      readAddr2_xhdl350 := "00000000000000";    
      readAddr3_xhdl351 := "00000000000000";    
      readAddr4_xhdl352 := "00000000000000";    
      readAddr5_xhdl353 := "00000000000000";    
      readAddr6_xhdl354 := "00000000000000";    
      readAddr7_xhdl355 := "00000000000000";    
      readAddr8_xhdl356 := "00000000000000";    
      readAddr9_xhdl357 := "00000000000000";    
      readAddr10_xhdl358 := "00000000000000";    
      readAddr11_xhdl359 := "00000000000000";    
      readAddr12_xhdl360 := "00000000000000";    
      readAddr13_xhdl361 := "00000000000000";    
      readAddr14_xhdl362 := "00000000000000";    
      readAddr15_xhdl363 := "00000000000000";    
      readAddr16_xhdl364 := "00000000000000";    
      readAddr17_xhdl365 := "00000000000000";    
      readAddr18_xhdl366 := "00000000000000";    
      readAddr19_xhdl367 := "00000000000000";    
      readAddr20_xhdl368 := "00000000000000";    
      readAddr21_xhdl369 := "00000000000000";    
      readAddr22_xhdl370 := "00000000000000";    
      readAddr23_xhdl371 := "00000000000000";    
      readAddr24_xhdl372 := "00000000000000";    
      readAddr25_xhdl373 := "00000000000000";    
      readAddr26_xhdl374 := "00000000000000";    
      readAddr27_xhdl375 := "00000000000000";    
      readAddr28_xhdl376 := "00000000000000";    
      readAddr29_xhdl377 := "00000000000000";    
      readAddr30_xhdl378 := "00000000000000";    
      readAddr31_xhdl379 := "00000000000000";    
      readAddr32_xhdl380 := "00000000000000";    
      readAddr33_xhdl381 := "00000000000000";    
      readAddr34_xhdl382 := "00000000000000";    
      readAddr35_xhdl383 := "00000000000000";    
      readAddr36_xhdl384 := "00000000000000";    
      readAddr37_xhdl385 := "00000000000000";    
      readAddr38_xhdl386 := "00000000000000";    
      readAddr39_xhdl387 := "00000000000000";    
      readAddr40_xhdl388 := "00000000000000";    
      readAddr41_xhdl389 := "00000000000000";    
      readAddr42_xhdl390 := "00000000000000";    
      readAddr43_xhdl391 := "00000000000000";    
      readAddr44_xhdl392 := "00000000000000";    
      readAddr45_xhdl393 := "00000000000000";    
      readAddr46_xhdl394 := "00000000000000";    
      readAddr47_xhdl395 := "00000000000000";    
      readAddr48_xhdl396 := "00000000000000";    
      readAddr49_xhdl397 := "00000000000000";    
      readAddr50_xhdl398 := "00000000000000";    
      readAddr51_xhdl399 := "00000000000000";    
      readAddr52_xhdl400 := "00000000000000";    
      readAddr53_xhdl401 := "00000000000000";    
      readAddr54_xhdl402 := "00000000000000";    
      readAddr55_xhdl403 := "00000000000000";    
      readAddr56_xhdl404 := "00000000000000";    
      readAddr57_xhdl405 := "00000000000000";    
      readAddr58_xhdl406 := "00000000000000";    
      readAddr59_xhdl407 := "00000000000000";    
      readAddr60_xhdl408 := "00000000000000";    
      readAddr61_xhdl409 := "00000000000000";    
      readAddr62_xhdl410 := "00000000000000";    
      readAddr63_xhdl411 := "00000000000000";    
      readAddr64_xhdl412 := "00000000000000";    
      readAddr65_xhdl413 := "00000000000000";    
      readAddr66_xhdl414 := "00000000000000";    
      readAddr67_xhdl415 := "00000000000000";    
      readAddr68_xhdl416 := "00000000000000";    
      readData_xhdl1_xhdl417 := (OTHERS => '0');    
      CASE DEPTH IS
         WHEN 2048 =>
                  width1_xhdl4 := "011";    
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  wen_a1_xhdl73 := '0' & wen;    
                  readData_xhdl1_xhdl417 := readData1(7 DOWNTO 0);    
         WHEN 4096 =>
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "0000" |
                          "0001" =>
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN "0010" |
                          "0011" =>
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN OTHERS  =>
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:12])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (ckRdAddr[13:12])               
                  
                  
         WHEN 6144 =>
                  width2_xhdl5 := "011";    
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr2_xhdl281 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr2_xhdl350 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData2_xhdl212 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "0000" |
                          "0001" =>
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN "0010" |
                          "0011" =>
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100" |
                          "0101" =>
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN OTHERS  =>
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:12])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN "0100" |
                          "0101" =>
                              readData_xhdl1_xhdl417 := readData2(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:12])
                  
                  
         WHEN 8192 =>
                  width3_xhdl6 := "011";    
                  width2_xhdl5 := "011";    
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr3_xhdl282 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr2_xhdl281 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr3_xhdl351 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr2_xhdl350 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData3_xhdl213 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData2_xhdl212 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "0110" |
                          "0111" =>
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100" |
                          "0101" =>
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010" |
                          "0011" =>
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000" |
                          "0001" =>
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:12])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "0110" |
                          "0111" =>
                              readData_xhdl1_xhdl417 := readData3(7 
                              DOWNTO 0);    
                     WHEN "0100" |
                          "0101" =>
                              readData_xhdl1_xhdl417 := readData2(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:12])
                  
                  
         WHEN 10240 =>
                  width4_xhdl7 := "011";    
                  width3_xhdl6 := "011";    
                  width2_xhdl5 := "011";    
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr4_xhdl283 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr3_xhdl282 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr2_xhdl281 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr4_xhdl352 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr3_xhdl351 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr2_xhdl350 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData4_xhdl214 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData3_xhdl213 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData2_xhdl212 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "1000" |
                          "1001" =>
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110" |
                          "0111" =>
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100" |
                          "0101" =>
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010" |
                          "0011" =>
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000" |
                          "0001" =>
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "1000" |
                          "1001" =>
                              readData_xhdl1_xhdl417 := readData4(7 
                              DOWNTO 0);    
                     WHEN "0110" |
                          "0111" =>
                              readData_xhdl1_xhdl417 := readData3(7 
                              DOWNTO 0);    
                     WHEN "0100" |
                          "0101" =>
                              readData_xhdl1_xhdl417 := readData2(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  
         WHEN 12288 =>
                  width5_xhdl8 := "011";    
                  width4_xhdl7 := "011";    
                  width3_xhdl6 := "011";    
                  width2_xhdl5 := "011";    
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr5_xhdl284 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr4_xhdl283 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr3_xhdl282 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr2_xhdl281 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr5_xhdl353 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr4_xhdl352 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr3_xhdl351 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr2_xhdl350 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData5_xhdl215 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData4_xhdl214 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData3_xhdl213 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData2_xhdl212 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "1010" |
                          "1011" =>
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000" |
                          "1001" =>
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110" |
                          "0111" =>
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100" |
                          "0101" =>
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010" |
                          "0011" =>
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000" |
                          "0001" =>
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "1010" |
                          "1011" =>
                              readData_xhdl1_xhdl417 := readData5(7 
                              DOWNTO 0);    
                     WHEN "1000" |
                          "1001" =>
                              readData_xhdl1_xhdl417 := readData4(7 
                              DOWNTO 0);    
                     WHEN "0110" |
                          "0111" =>
                              readData_xhdl1_xhdl417 := readData3(7 
                              DOWNTO 0);    
                     WHEN "0100" |
                          "0101" =>
                              readData_xhdl1_xhdl417 := readData2(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  
         WHEN 14336 =>
                  width6_xhdl9 := "011";    
                  width5_xhdl8 := "011";    
                  width4_xhdl7 := "011";    
                  width3_xhdl6 := "011";    
                  width2_xhdl5 := "011";    
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr6_xhdl285 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr5_xhdl284 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr4_xhdl283 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr3_xhdl282 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr2_xhdl281 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr6_xhdl354 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr5_xhdl353 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr4_xhdl352 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr3_xhdl351 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr2_xhdl350 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData6_xhdl216 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData5_xhdl215 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData4_xhdl214 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData3_xhdl213 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData2_xhdl212 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "1100" |
                          "1101" =>
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010" |
                          "1011" =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000" |
                          "1001" =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110" |
                          "0111" =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100" |
                          "0101" =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010" |
                          "0011" =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000" |
                          "0001" =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "1100" |
                          "1101" =>
                              readData_xhdl1_xhdl417 := readData6(7 
                              DOWNTO 0);    
                     WHEN "1010" |
                          "1011" =>
                              readData_xhdl1_xhdl417 := readData5(7 
                              DOWNTO 0);    
                     WHEN "1000" |
                          "1001" =>
                              readData_xhdl1_xhdl417 := readData4(7 
                              DOWNTO 0);    
                     WHEN "0110" |
                          "0111" =>
                              readData_xhdl1_xhdl417 := readData3(7 
                              DOWNTO 0);    
                     WHEN "0100" |
                          "0101" =>
                              readData_xhdl1_xhdl417 := readData2(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  
         WHEN 16384 =>
                  width7_xhdl10 := "011";    
                  width6_xhdl9 := "011";    
                  width5_xhdl8 := "011";    
                  width4_xhdl7 := "011";    
                  width3_xhdl6 := "011";    
                  width2_xhdl5 := "011";    
                  width1_xhdl4 := "011";    
                  width0_xhdl3 := "011";    
                  writeAddr7_xhdl286 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr6_xhdl285 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr5_xhdl284 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr4_xhdl283 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr3_xhdl282 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr2_xhdl281 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr1_xhdl280 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr0_xhdl279 := writeAddr(10 DOWNTO 0) & "000";  
                  readAddr7_xhdl355 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr6_xhdl354 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr5_xhdl353 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr4_xhdl352 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr3_xhdl351 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr2_xhdl350 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr1_xhdl349 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr0_xhdl348 := readAddr(10 DOWNTO 0) & "000";    
                  writeData7_xhdl217 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData6_xhdl216 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData5_xhdl215 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData4_xhdl214 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData3_xhdl213 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData2_xhdl212 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData1_xhdl211 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData0_xhdl210 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  CASE writeAddr(13 DOWNTO 10) IS
                     WHEN "1110" |
                          "1111" =>
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100" |
                          "1101" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010" |
                          "1011" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000" |
                          "1001" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110" |
                          "0111" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100" |
                          "0101" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010" |
                          "0011" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000" |
                          "0001" =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  CASE ckRdAddr(13 DOWNTO 10) IS
                     WHEN "1110" |
                          "1111" =>
                              readData_xhdl1_xhdl417 := readData7(7 
                              DOWNTO 0);    
                     WHEN "1100" |
                          "1101" =>
                              readData_xhdl1_xhdl417 := readData6(7 
                              DOWNTO 0);    
                     WHEN "1010" |
                          "1011" =>
                              readData_xhdl1_xhdl417 := readData5(7 
                              DOWNTO 0);    
                     WHEN "1000" |
                          "1001" =>
                              readData_xhdl1_xhdl417 := readData4(7 
                              DOWNTO 0);    
                     WHEN "0110" |
                          "0111" =>
                              readData_xhdl1_xhdl417 := readData3(7 
                              DOWNTO 0);    
                     WHEN "0100" |
                          "0101" =>
                              readData_xhdl1_xhdl417 := readData2(7 
                              DOWNTO 0);    
                     WHEN "0010" |
                          "0011" =>
                              readData_xhdl1_xhdl417 := readData1(7 
                              DOWNTO 0);    
                     WHEN "0000" |
                          "0001" =>
                              readData_xhdl1_xhdl417 := readData0(7 
                              DOWNTO 0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  
         WHEN 18432 =>
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "10000" |
                          "10001" =>
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  
         WHEN 20480 =>
                  width9_xhdl12 := "011";    
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr9_xhdl288 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData9_xhdl219 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "10010" |
                          "10011" =>
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000" |
                          "10001" =>
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "10010" |
                          "10011" =>
                              readData_xhdl1_xhdl417 := readData9(7 
                              DOWNTO 0);    
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[13:10])
                  
                  
         WHEN 22528 =>
                  width10_xhdl13 := "011";    
                  width9_xhdl12 := "011";    
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr10_xhdl289 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr9_xhdl288 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr9_xhdl357 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData10_xhdl220 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData9_xhdl219 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "10100" |
                          "10101" =>
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10010" |
                          "10011" =>
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000" |
                          "10001" =>
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "10100" |
                          "10101" =>
                              readData_xhdl1_xhdl417 := readData10(7 
                              DOWNTO 0);    
                     WHEN "10010" |
                          "10011" =>
                              readData_xhdl1_xhdl417 := readData9(7 
                              DOWNTO 0);    
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
         WHEN 24576 =>
                  width11_xhdl14 := "011";    
                  width10_xhdl13 := "011";    
                  width9_xhdl12 := "011";    
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr11_xhdl290 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr10_xhdl289 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr9_xhdl288 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr10_xhdl358 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr9_xhdl357 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData11_xhdl221 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData10_xhdl220 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData9_xhdl219 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "10110" |
                          "10111" =>
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10100" |
                          "10101" =>
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10010" |
                          "10011" =>
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000" |
                          "10001" =>
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "10110" |
                          "10111" =>
                              readData_xhdl1_xhdl417 := readData11(7 
                              DOWNTO 0);    
                     WHEN "10100" |
                          "10101" =>
                              readData_xhdl1_xhdl417 := readData10(7 
                              DOWNTO 0);    
                     WHEN "10010" |
                          "10011" =>
                              readData_xhdl1_xhdl417 := readData9(7 
                              DOWNTO 0);    
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
         WHEN 26624 =>
                  width12_xhdl15 := "011";    
                  width11_xhdl14 := "011";    
                  width10_xhdl13 := "011";    
                  width9_xhdl12 := "011";    
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr12_xhdl291 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr11_xhdl290 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr10_xhdl289 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr9_xhdl288 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr11_xhdl359 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr10_xhdl358 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr9_xhdl357 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData12_xhdl222 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData11_xhdl221 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData10_xhdl220 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData9_xhdl219 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "11000" |
                          "11001" =>
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10110" |
                          "10111" =>
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10100" |
                          "10101" =>
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10010" |
                          "10011" =>
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000" |
                          "10001" =>
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "11000" |
                          "11001" =>
                              readData_xhdl1_xhdl417 := readData12(7 
                              DOWNTO 0);    
                     WHEN "10110" |
                          "10111" =>
                              readData_xhdl1_xhdl417 := readData11(7 
                              DOWNTO 0);    
                     WHEN "10100" |
                          "10101" =>
                              readData_xhdl1_xhdl417 := readData10(7 
                              DOWNTO 0);    
                     WHEN "10010" |
                          "10011" =>
                              readData_xhdl1_xhdl417 := readData9(7 
                              DOWNTO 0);    
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
         WHEN 28672 =>
                  width13_xhdl16 := "011";    
                  width12_xhdl15 := "011";    
                  width11_xhdl14 := "011";    
                  width10_xhdl13 := "011";    
                  width9_xhdl12 := "011";    
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr13_xhdl292 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr12_xhdl291 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr11_xhdl290 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr10_xhdl289 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr9_xhdl288 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr12_xhdl360 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr11_xhdl359 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr10_xhdl358 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr9_xhdl357 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData13_xhdl223 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData12_xhdl222 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData11_xhdl221 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData10_xhdl220 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData9_xhdl219 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "11010" |
                          "11011" =>
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "11000" |
                          "11001" =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10110" |
                          "10111" =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10100" |
                          "10101" =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10010" |
                          "10011" =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000" |
                          "10001" =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "11010" |
                          "11011" =>
                              readData_xhdl1_xhdl417 := readData13(7 
                              DOWNTO 0);    
                     WHEN "11000" |
                          "11001" =>
                              readData_xhdl1_xhdl417 := readData12(7 
                              DOWNTO 0);    
                     WHEN "10110" |
                          "10111" =>
                              readData_xhdl1_xhdl417 := readData11(7 
                              DOWNTO 0);    
                     WHEN "10100" |
                          "10101" =>
                              readData_xhdl1_xhdl417 := readData10(7 
                              DOWNTO 0);    
                     WHEN "10010" |
                          "10011" =>
                              readData_xhdl1_xhdl417 := readData9(7 
                              DOWNTO 0);    
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
         WHEN 30720 =>
                  width14_xhdl17 := "011";    
                  width13_xhdl16 := "011";    
                  width12_xhdl15 := "011";    
                  width11_xhdl14 := "011";    
                  width10_xhdl13 := "011";    
                  width9_xhdl12 := "011";    
                  width8_xhdl11 := "011";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr14_xhdl293 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr13_xhdl292 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr12_xhdl291 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr11_xhdl290 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr10_xhdl289 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr9_xhdl288 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr8_xhdl287 := writeAddr(10 DOWNTO 0) & "000";  
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr13_xhdl361 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr12_xhdl360 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr11_xhdl359 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr10_xhdl358 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr9_xhdl357 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr8_xhdl356 := readAddr(10 DOWNTO 0) & "000";    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData14_xhdl224 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData13_xhdl223 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData12_xhdl222 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData11_xhdl221 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData10_xhdl220 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData9_xhdl219 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData8_xhdl218 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "11100" |
                          "11101" =>
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "11010" |
                          "11011" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "11000" |
                          "11001" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10110" |
                          "10111" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10100" |
                          "10101" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10010" |
                          "10011" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000" |
                          "10001" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "11100" |
                          "11101" =>
                              readData_xhdl1_xhdl417 := readData14(7 
                              DOWNTO 0);    
                     WHEN "11010" |
                          "11011" =>
                              readData_xhdl1_xhdl417 := readData13(7 
                              DOWNTO 0);    
                     WHEN "11000" |
                          "11001" =>
                              readData_xhdl1_xhdl417 := readData12(7 
                              DOWNTO 0);    
                     WHEN "10110" |
                          "10111" =>
                              readData_xhdl1_xhdl417 := readData11(7 
                              DOWNTO 0);    
                     WHEN "10100" |
                          "10101" =>
                              readData_xhdl1_xhdl417 := readData10(7 
                              DOWNTO 0);    
                     WHEN "10010" |
                          "10011" =>
                              readData_xhdl1_xhdl417 := readData9(7 
                              DOWNTO 0);    
                     WHEN "10000" |
                          "10001" =>
                              readData_xhdl1_xhdl417 := readData8(7 
                              DOWNTO 0);    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
         WHEN 32768 =>
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(14 DOWNTO 10) IS
                     WHEN "10000" |
                          "10001" |
                          "10010" |
                          "10011" |
                          "10100" |
                          "10101" |
                          "10110" |
                          "10111" |
                          "11000" |
                          "11001" |
                          "11010" |
                          "11011" |
                          "11100" |
                          "11101" |
                          "11110" |
                          "11111" =>
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(14 DOWNTO 10) IS
                     WHEN "10000" |
                          "10001" |
                          "10010" |
                          "10011" |
                          "10100" |
                          "10101" |
                          "10110" |
                          "10111" |
                          "11000" |
                          "11001" |
                          "11010" |
                          "11011" |
                          "11100" |
                          "11101" |
                          "11110" |
                          "11111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "00000" |
                          "00001" |
                          "00010" |
                          "00011" |
                          "00100" |
                          "00101" |
                          "00110" |
                          "00111" |
                          "01000" |
                          "01001" |
                          "01010" |
                          "01011" |
                          "01100" |
                          "01101" |
                          "01110" |
                          "01111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
          
                  
         WHEN 34816 =>
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "100000" |
                          "100001" =>
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[14:10])
                  
                  
         WHEN 36864 =>
                  width17_xhdl20 := "011";    
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr17_xhdl296 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData17_xhdl227 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "100010" |
                          "100011" =>
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" =>
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "100010" |
                          "100011" =>
                              readData_xhdl1_xhdl417 := readData17(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 38912 =>
                  width18_xhdl21 := "011";    
                  width17_xhdl20 := "011";    
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr18_xhdl297 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr17_xhdl296 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr17_xhdl365 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData18_xhdl228 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData17_xhdl227 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "100100" |
                          "100101" =>
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100010" |
                          "100011" =>
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" =>
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "100100" |
                          "100101" =>
                              readData_xhdl1_xhdl417 := readData18(7 
                              DOWNTO 0);    
                     WHEN "100010" |
                          "100011" =>
                              readData_xhdl1_xhdl417 := readData17(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 40960 =>
                  width19_xhdl22 := "011";    
                  width18_xhdl21 := "011";    
                  width17_xhdl20 := "011";    
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr19_xhdl298 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr18_xhdl297 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr17_xhdl296 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr18_xhdl366 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr17_xhdl365 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData19_xhdl229 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData18_xhdl228 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData17_xhdl227 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "100110" |
                          "100111" =>
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100100" |
                          "100101" =>
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100010" |
                          "100011" =>
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" =>
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "100110" |
                          "100111" =>
                              readData_xhdl1_xhdl417 := readData19(7 
                              DOWNTO 0);    
                     WHEN "100100" |
                          "100101" =>
                              readData_xhdl1_xhdl417 := readData18(7 
                              DOWNTO 0);    
                     WHEN "100010" |
                          "100011" =>
                              readData_xhdl1_xhdl417 := readData17(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 43008 =>
                  width20_xhdl23 := "011";    
                  width19_xhdl22 := "011";    
                  width18_xhdl21 := "011";    
                  width17_xhdl20 := "011";    
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr20_xhdl299 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr19_xhdl298 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr18_xhdl297 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr17_xhdl296 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr19_xhdl367 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr18_xhdl366 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr17_xhdl365 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData20_xhdl230 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData19_xhdl229 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData18_xhdl228 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData17_xhdl227 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "101000" |
                          "101001" =>
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100110" |
                          "100111" =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100100" |
                          "100101" =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100010" |
                          "100011" =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "101000" |
                          "101001" =>
                              readData_xhdl1_xhdl417 := readData20(7 
                              DOWNTO 0);    
                     WHEN "100110" |
                          "100111" =>
                              readData_xhdl1_xhdl417 := readData19(7 
                              DOWNTO 0);    
                     WHEN "100100" |
                          "100101" =>
                              readData_xhdl1_xhdl417 := readData18(7 
                              DOWNTO 0);    
                     WHEN "100010" |
                          "100011" =>
                              readData_xhdl1_xhdl417 := readData17(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 45056 =>
                  width21_xhdl24 := "011";    
                  width20_xhdl23 := "011";    
                  width19_xhdl22 := "011";    
                  width18_xhdl21 := "011";    
                  width17_xhdl20 := "011";    
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr21_xhdl300 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr20_xhdl299 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr19_xhdl298 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr18_xhdl297 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr17_xhdl296 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr20_xhdl368 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr19_xhdl367 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr18_xhdl366 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr17_xhdl365 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData21_xhdl231 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData20_xhdl230 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData19_xhdl229 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData18_xhdl228 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData17_xhdl227 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "101010" |
                          "101011" =>
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "101000" |
                          "101001" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100110" |
                          "100111" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100100" |
                          "100101" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100010" |
                          "100011" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "101010" |
                          "101011" =>
                              readData_xhdl1_xhdl417 := readData21(7 
                              DOWNTO 0);    
                     WHEN "101000" |
                          "101001" =>
                              readData_xhdl1_xhdl417 := readData20(7 
                              DOWNTO 0);    
                     WHEN "100110" |
                          "100111" =>
                              readData_xhdl1_xhdl417 := readData19(7 
                              DOWNTO 0);    
                     WHEN "100100" |
                          "100101" =>
                              readData_xhdl1_xhdl417 := readData18(7 
                              DOWNTO 0);    
                     WHEN "100010" |
                          "100011" =>
                              readData_xhdl1_xhdl417 := readData17(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 47104 =>
                  width22_xhdl25 := "011";    
                  width21_xhdl24 := "011";    
                  width20_xhdl23 := "011";    
                  width19_xhdl22 := "011";    
                  width18_xhdl21 := "011";    
                  width17_xhdl20 := "011";    
                  width16_xhdl19 := "011";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr22_xhdl301 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr21_xhdl300 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr20_xhdl299 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr19_xhdl298 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr18_xhdl297 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr17_xhdl296 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr16_xhdl295 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr21_xhdl369 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr20_xhdl368 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr19_xhdl367 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr18_xhdl366 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr17_xhdl365 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr16_xhdl364 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData22_xhdl232 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData21_xhdl231 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData20_xhdl230 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData19_xhdl229 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData18_xhdl228 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData17_xhdl227 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData16_xhdl226 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "101100" |
                          "101101" =>
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "101010" |
                          "101011" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "101000" |
                          "101001" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100110" |
                          "100111" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100100" |
                          "100101" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100010" |
                          "100011" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "101100" |
                          "101101" =>
                              readData_xhdl1_xhdl417 := readData22(7 
                              DOWNTO 0);    
                     WHEN "101010" |
                          "101011" =>
                              readData_xhdl1_xhdl417 := readData21(7 
                              DOWNTO 0);    
                     WHEN "101000" |
                          "101001" =>
                              readData_xhdl1_xhdl417 := readData20(7 
                              DOWNTO 0);    
                     WHEN "100110" |
                          "100111" =>
                              readData_xhdl1_xhdl417 := readData19(7 
                              DOWNTO 0);    
                     WHEN "100100" |
                          "100101" =>
                              readData_xhdl1_xhdl417 := readData18(7 
                              DOWNTO 0);    
                     WHEN "100010" |
                          "100011" =>
                              readData_xhdl1_xhdl417 := readData17(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" =>
                              readData_xhdl1_xhdl417 := readData16(7 
                              DOWNTO 0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 49152 =>
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 51200 =>
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "110000" |
                          "110001" =>
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 53248 =>
                  width25_xhdl28 := "011";    
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr25_xhdl304 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData25_xhdl235 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "110010" |
                          "110011" =>
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110000" |
                          "110001" =>
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "110010" |
                          "110011" =>
                              readData_xhdl1_xhdl417 := readData25(7 
                              DOWNTO 0);    
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 55296 =>
                  width26_xhdl29 := "011";    
                  width25_xhdl28 := "011";    
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr26_xhdl305 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr25_xhdl304 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr25_xhdl373 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData26_xhdl236 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData25_xhdl235 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "110100" |
                          "110101" =>
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110010" |
                          "110011" =>
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110000" |
                          "110001" =>
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "110100" |
                          "110101" =>
                              readData_xhdl1_xhdl417 := readData26(7 
                              DOWNTO 0);    
                     WHEN "110010" |
                          "110011" =>
                              readData_xhdl1_xhdl417 := readData25(7 
                              DOWNTO 0);    
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 57344 =>
                  width27_xhdl30 := "011";    
                  width26_xhdl29 := "011";    
                  width25_xhdl28 := "011";    
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr27_xhdl306 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr26_xhdl305 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr25_xhdl304 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr26_xhdl374 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr25_xhdl373 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData27_xhdl237 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData26_xhdl236 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData25_xhdl235 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "110110" |
                          "110111" =>
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110100" |
                          "110101" =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110010" |
                          "110011" =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110000" |
                          "110001" =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "110110" |
                          "110111" =>
                              readData_xhdl1_xhdl417 := readData27(7 
                              DOWNTO 0);    
                     WHEN "110100" |
                          "110101" =>
                              readData_xhdl1_xhdl417 := readData26(7 
                              DOWNTO 0);    
                     WHEN "110010" |
                          "110011" =>
                              readData_xhdl1_xhdl417 := readData25(7 
                              DOWNTO 0);    
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 59392 =>
                  width28_xhdl31 := "011";    
                  width27_xhdl30 := "011";    
                  width26_xhdl29 := "011";    
                  width25_xhdl28 := "011";    
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr28_xhdl307 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr27_xhdl306 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr26_xhdl305 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr25_xhdl304 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr27_xhdl375 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr26_xhdl374 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr25_xhdl373 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData28_xhdl238 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData27_xhdl237 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData26_xhdl236 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData25_xhdl235 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "111000" |
                          "111001" =>
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110110" |
                          "110111" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110100" |
                          "110101" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110010" |
                          "110011" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110000" |
                          "110001" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "111000" |
                          "111001" =>
                              readData_xhdl1_xhdl417 := readData28(7 
                              DOWNTO 0);    
                     WHEN "110110" |
                          "110111" =>
                              readData_xhdl1_xhdl417 := readData27(7 
                              DOWNTO 0);    
                     WHEN "110100" |
                          "110101" =>
                              readData_xhdl1_xhdl417 := readData26(7 
                              DOWNTO 0);    
                     WHEN "110010" |
                          "110011" =>
                              readData_xhdl1_xhdl417 := readData25(7 
                              DOWNTO 0);    
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 61440 =>
                  width29_xhdl32 := "011";    
                  width28_xhdl31 := "011";    
                  width27_xhdl30 := "011";    
                  width26_xhdl29 := "011";    
                  width25_xhdl28 := "011";    
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr29_xhdl308 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr28_xhdl307 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr27_xhdl306 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr26_xhdl305 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr25_xhdl304 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr28_xhdl376 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr27_xhdl375 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr26_xhdl374 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr25_xhdl373 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData29_xhdl239 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData28_xhdl238 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData27_xhdl237 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData26_xhdl236 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData25_xhdl235 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "111010" |
                          "111011" =>
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "111000" |
                          "111001" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110110" |
                          "110111" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110100" |
                          "110101" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110010" |
                          "110011" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110000" |
                          "110001" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "111010" |
                          "111011" =>
                              readData_xhdl1_xhdl417 := readData29(7 
                              DOWNTO 0);    
                     WHEN "111000" |
                          "111001" =>
                              readData_xhdl1_xhdl417 := readData28(7 
                              DOWNTO 0);    
                     WHEN "110110" |
                          "110111" =>
                              readData_xhdl1_xhdl417 := readData27(7 
                              DOWNTO 0);    
                     WHEN "110100" |
                          "110101" =>
                              readData_xhdl1_xhdl417 := readData26(7 
                              DOWNTO 0);    
                     WHEN "110010" |
                          "110011" =>
                              readData_xhdl1_xhdl417 := readData25(7 
                              DOWNTO 0);    
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 63488 =>
                  width30_xhdl33 := "011";    
                  width29_xhdl32 := "011";    
                  width28_xhdl31 := "011";    
                  width27_xhdl30 := "011";    
                  width26_xhdl29 := "011";    
                  width25_xhdl28 := "011";    
                  width24_xhdl27 := "011";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr30_xhdl309 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr29_xhdl308 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr28_xhdl307 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr27_xhdl306 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr26_xhdl305 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr25_xhdl304 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr24_xhdl303 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr29_xhdl377 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr28_xhdl376 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr27_xhdl375 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr26_xhdl374 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr25_xhdl373 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr24_xhdl372 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData30_xhdl240 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData29_xhdl239 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData28_xhdl238 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData27_xhdl237 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData26_xhdl236 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData25_xhdl235 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData24_xhdl234 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "111100" |
                          "111101" =>
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "111010" |
                          "111011" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "111000" |
                          "111001" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110110" |
                          "110111" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110100" |
                          "110101" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110010" |
                          "110011" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "110000" |
                          "110001" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "111100" |
                          "111101" =>
                              readData_xhdl1_xhdl417 := readData30(7 
                              DOWNTO 0);    
                     WHEN "111010" |
                          "111011" =>
                              readData_xhdl1_xhdl417 := readData29(7 
                              DOWNTO 0);    
                     WHEN "111000" |
                          "111001" =>
                              readData_xhdl1_xhdl417 := readData28(7 
                              DOWNTO 0);    
                     WHEN "110110" |
                          "110111" =>
                              readData_xhdl1_xhdl417 := readData27(7 
                              DOWNTO 0);    
                     WHEN "110100" |
                          "110101" =>
                              readData_xhdl1_xhdl417 := readData26(7 
                              DOWNTO 0);    
                     WHEN "110010" |
                          "110011" =>
                              readData_xhdl1_xhdl417 := readData25(7 
                              DOWNTO 0);    
                     WHEN "110000" |
                          "110001" =>
                              readData_xhdl1_xhdl417 := readData24(7 
                              DOWNTO 0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 65536 =>
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(15 DOWNTO 10) IS
                     WHEN "110000" |
                          "110001" |
                          "110010" |
                          "110011" |
                          "110100" |
                          "110101" |
                          "110110" |
                          "110111" |
                          "111000" |
                          "111001" |
                          "111010" |
                          "111011" |
                          "111100" |
                          "111101" |
                          "111110" |
                          "111111" =>
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  CASE ckRdAddr(15 DOWNTO 10) IS
                     WHEN "110000" |
                          "110001" |
                          "110010" |
                          "110011" |
                          "110100" |
                          "110101" |
                          "110110" |
                          "110111" |
                          "111000" |
                          "111001" |
                          "111010" |
                          "111011" |
                          "111100" |
                          "111101" |
                          "111110" |
                          "111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "100000" |
                          "100001" |
                          "100010" |
                          "100011" |
                          "100100" |
                          "100101" |
                          "100110" |
                          "100111" |
                          "101000" |
                          "101001" |
                          "101010" |
                          "101011" |
                          "101100" |
                          "101101" |
                          "101110" |
                          "101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "010000" |
                          "010001" |
                          "010010" |
                          "010011" |
                          "010100" |
                          "010101" |
                          "010110" |
                          "010111" |
                          "011000" |
                          "011001" |
                          "011010" |
                          "011011" |
                          "011100" |
                          "011101" |
                          "011110" |
                          "011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "000000" |
                          "000001" |
                          "000010" |
                          "000011" |
                          "000100" |
                          "000101" |
                          "000110" |
                          "000111" |
                          "001000" |
                          "001001" |
                          "001010" |
                          "001011" |
                          "001100" |
                          "001101" |
                          "001110" |
                          "001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[15:10])
                  
                  
         WHEN 67584 =>
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 69632 =>
                  width33_xhdl36 := "011";    
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr33_xhdl312 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData33_xhdl243 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1000010" |
                          "1000011" =>
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1000010" |
                          "1000011" =>
                              readData_xhdl1_xhdl417 := readData33(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 71680 =>
                  width34_xhdl37 := "011";    
                  width33_xhdl36 := "011";    
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr34_xhdl313 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr33_xhdl312 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr33_xhdl381 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData34_xhdl244 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData33_xhdl243 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1000100" |
                          "1000101" =>
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000010" |
                          "1000011" =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1000100" |
                          "1000101" =>
                              readData_xhdl1_xhdl417 := readData34(7 
                              DOWNTO 0);    
                     WHEN "1000010" |
                          "1000011" =>
                              readData_xhdl1_xhdl417 := readData33(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 73728 =>
                  width35_xhdl38 := "011";    
                  width34_xhdl37 := "011";    
                  width33_xhdl36 := "011";    
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr35_xhdl314 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr34_xhdl313 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr33_xhdl312 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr34_xhdl382 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr33_xhdl381 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData35_xhdl245 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData34_xhdl244 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData33_xhdl243 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1000110" |
                          "1000111" =>
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000100" |
                          "1000101" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000010" |
                          "1000011" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1000110" |
                          "1000111" =>
                              readData_xhdl1_xhdl417 := readData35(7 
                              DOWNTO 0);    
                     WHEN "1000100" |
                          "1000101" =>
                              readData_xhdl1_xhdl417 := readData34(7 
                              DOWNTO 0);    
                     WHEN "1000010" |
                          "1000011" =>
                              readData_xhdl1_xhdl417 := readData33(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 75776 =>
                  width36_xhdl39 := "011";    
                  width35_xhdl38 := "011";    
                  width34_xhdl37 := "011";    
                  width33_xhdl36 := "011";    
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr36_xhdl315 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr35_xhdl314 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr34_xhdl313 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr33_xhdl312 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr35_xhdl383 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr34_xhdl382 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr33_xhdl381 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData36_xhdl246 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData35_xhdl245 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData34_xhdl244 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData33_xhdl243 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1001000" |
                          "1001001" =>
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000110" |
                          "1000111" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000100" |
                          "1000101" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000010" |
                          "1000011" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1001000" |
                          "1001001" =>
                              readData_xhdl1_xhdl417 := readData36(7 
                              DOWNTO 0);    
                     WHEN "1000110" |
                          "1000111" =>
                              readData_xhdl1_xhdl417 := readData35(7 
                              DOWNTO 0);    
                     WHEN "1000100" |
                          "1000101" =>
                              readData_xhdl1_xhdl417 := readData34(7 
                              DOWNTO 0);    
                     WHEN "1000010" |
                          "1000011" =>
                              readData_xhdl1_xhdl417 := readData33(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 77824 =>
                  width37_xhdl40 := "011";    
                  width36_xhdl39 := "011";    
                  width35_xhdl38 := "011";    
                  width34_xhdl37 := "011";    
                  width33_xhdl36 := "011";    
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr37_xhdl316 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr36_xhdl315 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr35_xhdl314 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr34_xhdl313 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr33_xhdl312 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr36_xhdl384 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr35_xhdl383 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr34_xhdl382 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr33_xhdl381 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData37_xhdl247 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData36_xhdl246 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData35_xhdl245 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData34_xhdl244 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData33_xhdl243 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1001010" |
                          "1001011" =>
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1001000" |
                          "1001001" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000110" |
                          "1000111" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000100" |
                          "1000101" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000010" |
                          "1000011" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1001010" |
                          "1001011" =>
                              readData_xhdl1_xhdl417 := readData37(7 
                              DOWNTO 0);    
                     WHEN "1001000" |
                          "1001001" =>
                              readData_xhdl1_xhdl417 := readData36(7 
                              DOWNTO 0);    
                     WHEN "1000110" |
                          "1000111" =>
                              readData_xhdl1_xhdl417 := readData35(7 
                              DOWNTO 0);    
                     WHEN "1000100" |
                          "1000101" =>
                              readData_xhdl1_xhdl417 := readData34(7 
                              DOWNTO 0);    
                     WHEN "1000010" |
                          "1000011" =>
                              readData_xhdl1_xhdl417 := readData33(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 79872 =>
                  width38_xhdl41 := "011";    
                  width37_xhdl40 := "011";    
                  width36_xhdl39 := "011";    
                  width35_xhdl38 := "011";    
                  width34_xhdl37 := "011";    
                  width33_xhdl36 := "011";    
                  width32_xhdl35 := "011";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr38_xhdl317 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr37_xhdl316 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr36_xhdl315 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr35_xhdl314 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr34_xhdl313 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr33_xhdl312 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr32_xhdl311 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr37_xhdl385 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr36_xhdl384 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr35_xhdl383 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr34_xhdl382 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr33_xhdl381 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr32_xhdl380 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData38_xhdl248 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData37_xhdl247 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData36_xhdl246 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData35_xhdl245 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData34_xhdl244 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData33_xhdl243 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData32_xhdl242 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1001100" |
                          "1001101" =>
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1001010" |
                          "1001011" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1001000" |
                          "1001001" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000110" |
                          "1000111" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000100" |
                          "1000101" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000010" |
                          "1000011" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1001100" |
                          "1001101" =>
                              readData_xhdl1_xhdl417 := readData38(7 
                              DOWNTO 0);    
                     WHEN "1001010" |
                          "1001011" =>
                              readData_xhdl1_xhdl417 := readData37(7 
                              DOWNTO 0);    
                     WHEN "1001000" |
                          "1001001" =>
                              readData_xhdl1_xhdl417 := readData36(7 
                              DOWNTO 0);    
                     WHEN "1000110" |
                          "1000111" =>
                              readData_xhdl1_xhdl417 := readData35(7 
                              DOWNTO 0);    
                     WHEN "1000100" |
                          "1000101" =>
                              readData_xhdl1_xhdl417 := readData34(7 
                              DOWNTO 0);    
                     WHEN "1000010" |
                          "1000011" =>
                              readData_xhdl1_xhdl417 := readData33(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" =>
                              readData_xhdl1_xhdl417 := readData32(7 
                              DOWNTO 0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 81920 =>
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 83968 =>
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 86016 =>
                  width41_xhdl44 := "011";    
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr41_xhdl320 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData41_xhdl251 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1010010" |
                          "1010011" =>
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1010010" |
                          "1010011" =>
                              readData_xhdl1_xhdl417 := readData41(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 88064 =>
                  width42_xhdl45 := "011";    
                  width41_xhdl44 := "011";    
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr42_xhdl321 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr41_xhdl320 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr41_xhdl389 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData42_xhdl252 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData41_xhdl251 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1010100" |
                          "1010101" =>
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010010" |
                          "1010011" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1010100" |
                          "1010101" =>
                              readData_xhdl1_xhdl417 := readData42(7 
                              DOWNTO 0);    
                     WHEN "1010010" |
                          "1010011" =>
                              readData_xhdl1_xhdl417 := readData41(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 90112 =>
                  width43_xhdl46 := "011";    
                  width42_xhdl45 := "011";    
                  width41_xhdl44 := "011";    
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr43_xhdl322 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr42_xhdl321 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr41_xhdl320 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr42_xhdl390 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr41_xhdl389 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData43_xhdl253 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData42_xhdl252 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData41_xhdl251 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1010110" |
                          "1010111" =>
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010100" |
                          "1010101" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010010" |
                          "1010011" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1010110" |
                          "1010111" =>
                              readData_xhdl1_xhdl417 := readData43(7 
                              DOWNTO 0);    
                     WHEN "1010100" |
                          "1010101" =>
                              readData_xhdl1_xhdl417 := readData42(7 
                              DOWNTO 0);    
                     WHEN "1010010" |
                          "1010011" =>
                              readData_xhdl1_xhdl417 := readData41(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 92160 =>
                  width44_xhdl47 := "011";    
                  width43_xhdl46 := "011";    
                  width42_xhdl45 := "011";    
                  width41_xhdl44 := "011";    
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr44_xhdl323 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr43_xhdl322 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr42_xhdl321 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr41_xhdl320 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr43_xhdl391 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr42_xhdl390 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr41_xhdl389 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData44_xhdl254 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData43_xhdl253 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData42_xhdl252 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData41_xhdl251 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1011000" |
                          "1011001" =>
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010110" |
                          "1010111" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010100" |
                          "1010101" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010010" |
                          "1010011" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1011000" |
                          "1011001" =>
                              readData_xhdl1_xhdl417 := readData44(7 
                              DOWNTO 0);    
                     WHEN "1010110" |
                          "1010111" =>
                              readData_xhdl1_xhdl417 := readData43(7 
                              DOWNTO 0);    
                     WHEN "1010100" |
                          "1010101" =>
                              readData_xhdl1_xhdl417 := readData42(7 
                              DOWNTO 0);    
                     WHEN "1010010" |
                          "1010011" =>
                              readData_xhdl1_xhdl417 := readData41(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 94208 =>
                  width45_xhdl48 := "011";    
                  width44_xhdl47 := "011";    
                  width43_xhdl46 := "011";    
                  width42_xhdl45 := "011";    
                  width41_xhdl44 := "011";    
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr45_xhdl324 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr44_xhdl323 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr43_xhdl322 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr42_xhdl321 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr41_xhdl320 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr44_xhdl392 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr43_xhdl391 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr42_xhdl390 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr41_xhdl389 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData45_xhdl255 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData44_xhdl254 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData43_xhdl253 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData42_xhdl252 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData41_xhdl251 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1011010" |
                          "1011011" =>
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1011000" |
                          "1011001" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010110" |
                          "1010111" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010100" |
                          "1010101" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010010" |
                          "1010011" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1011010" |
                          "1011011" =>
                              readData_xhdl1_xhdl417 := readData45(7 
                              DOWNTO 0);    
                     WHEN "1011000" |
                          "1011001" =>
                              readData_xhdl1_xhdl417 := readData44(7 
                              DOWNTO 0);    
                     WHEN "1010110" |
                          "1010111" =>
                              readData_xhdl1_xhdl417 := readData43(7 
                              DOWNTO 0);    
                     WHEN "1010100" |
                          "1010101" =>
                              readData_xhdl1_xhdl417 := readData42(7 
                              DOWNTO 0);    
                     WHEN "1010010" |
                          "1010011" =>
                              readData_xhdl1_xhdl417 := readData41(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 96256 =>
                  width46_xhdl49 := "011";    
                  width45_xhdl48 := "011";    
                  width44_xhdl47 := "011";    
                  width43_xhdl46 := "011";    
                  width42_xhdl45 := "011";    
                  width41_xhdl44 := "011";    
                  width40_xhdl43 := "011";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr46_xhdl325 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr45_xhdl324 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr44_xhdl323 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr43_xhdl322 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr42_xhdl321 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr41_xhdl320 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr40_xhdl319 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr45_xhdl393 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr44_xhdl392 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr43_xhdl391 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr42_xhdl390 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr41_xhdl389 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr40_xhdl388 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData46_xhdl256 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData45_xhdl255 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData44_xhdl254 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData43_xhdl253 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData42_xhdl252 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData41_xhdl251 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData40_xhdl250 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1011100" |
                          "1011101" =>
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1011010" |
                          "1011011" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1011000" |
                          "1011001" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010110" |
                          "1010111" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010100" |
                          "1010101" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010010" |
                          "1010011" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1011100" |
                          "1011101" =>
                              readData_xhdl1_xhdl417 := readData46(7 
                              DOWNTO 0);    
                     WHEN "1011010" |
                          "1011011" =>
                              readData_xhdl1_xhdl417 := readData45(7 
                              DOWNTO 0);    
                     WHEN "1011000" |
                          "1011001" =>
                              readData_xhdl1_xhdl417 := readData44(7 
                              DOWNTO 0);    
                     WHEN "1010110" |
                          "1010111" =>
                              readData_xhdl1_xhdl417 := readData43(7 
                              DOWNTO 0);    
                     WHEN "1010100" |
                          "1010101" =>
                              readData_xhdl1_xhdl417 := readData42(7 
                              DOWNTO 0);    
                     WHEN "1010010" |
                          "1010011" =>
                              readData_xhdl1_xhdl417 := readData41(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" =>
                              readData_xhdl1_xhdl417 := readData40(7 
                              DOWNTO 0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 98304 =>
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 100352 =>
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 102400 =>
                  width49_xhdl52 := "011";    
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr49_xhdl328 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData49_xhdl259 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1100010" |
                          "1100011" =>
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1100010" |
                          "1100011" =>
                              readData_xhdl1_xhdl417 := readData49(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 104448 =>
                  width50_xhdl53 := "011";    
                  width49_xhdl52 := "011";    
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr50_xhdl329 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr49_xhdl328 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr49_xhdl397 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData50_xhdl260 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData49_xhdl259 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1100100" |
                          "1100101" =>
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100010" |
                          "1100011" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1100100" |
                          "1100101" =>
                              readData_xhdl1_xhdl417 := readData50(7 
                              DOWNTO 0);    
                     WHEN "1100010" |
                          "1100011" =>
                              readData_xhdl1_xhdl417 := readData49(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 106496 =>
                  width51_xhdl54 := "011";    
                  width50_xhdl53 := "011";    
                  width49_xhdl52 := "011";    
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr51_xhdl330 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr50_xhdl329 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr49_xhdl328 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr50_xhdl398 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr49_xhdl397 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData51_xhdl261 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData50_xhdl260 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData49_xhdl259 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1100110" |
                          "1100111" =>
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100100" |
                          "1100101" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100010" |
                          "1100011" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1100110" |
                          "1100111" =>
                              readData_xhdl1_xhdl417 := readData51(7 
                              DOWNTO 0);    
                     WHEN "1100100" |
                          "1100101" =>
                              readData_xhdl1_xhdl417 := readData50(7 
                              DOWNTO 0);    
                     WHEN "1100010" |
                          "1100011" =>
                              readData_xhdl1_xhdl417 := readData49(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 108544 =>
                  width52_xhdl55 := "011";    
                  width51_xhdl54 := "011";    
                  width50_xhdl53 := "011";    
                  width49_xhdl52 := "011";    
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr52_xhdl331 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr51_xhdl330 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr50_xhdl329 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr49_xhdl328 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr51_xhdl399 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr50_xhdl398 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr49_xhdl397 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData52_xhdl262 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData51_xhdl261 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData50_xhdl260 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData49_xhdl259 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1101000" |
                          "1101001" =>
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100110" |
                          "1100111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100100" |
                          "1100101" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100010" |
                          "1100011" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1101000" |
                          "1101001" =>
                              readData_xhdl1_xhdl417 := readData52(7 
                              DOWNTO 0);    
                     WHEN "1100110" |
                          "1100111" =>
                              readData_xhdl1_xhdl417 := readData51(7 
                              DOWNTO 0);    
                     WHEN "1100100" |
                          "1100101" =>
                              readData_xhdl1_xhdl417 := readData50(7 
                              DOWNTO 0);    
                     WHEN "1100010" |
                          "1100011" =>
                              readData_xhdl1_xhdl417 := readData49(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 110592 =>
                  width53_xhdl56 := "011";    
                  width52_xhdl55 := "011";    
                  width51_xhdl54 := "011";    
                  width50_xhdl53 := "011";    
                  width49_xhdl52 := "011";    
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr53_xhdl332 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr52_xhdl331 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr51_xhdl330 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr50_xhdl329 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr49_xhdl328 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr52_xhdl400 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr51_xhdl399 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr50_xhdl398 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr49_xhdl397 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData53_xhdl263 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData52_xhdl262 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData51_xhdl261 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData50_xhdl260 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData49_xhdl259 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1101010" |
                          "1101011" =>
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1101000" |
                          "1101001" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100110" |
                          "1100111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100100" |
                          "1100101" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100010" |
                          "1100011" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1101010" |
                          "1101011" =>
                              readData_xhdl1_xhdl417 := readData53(7 
                              DOWNTO 0);    
                     WHEN "1101000" |
                          "1101001" =>
                              readData_xhdl1_xhdl417 := readData52(7 
                              DOWNTO 0);    
                     WHEN "1100110" |
                          "1100111" =>
                              readData_xhdl1_xhdl417 := readData51(7 
                              DOWNTO 0);    
                     WHEN "1100100" |
                          "1100101" =>
                              readData_xhdl1_xhdl417 := readData50(7 
                              DOWNTO 0);    
                     WHEN "1100010" |
                          "1100011" =>
                              readData_xhdl1_xhdl417 := readData49(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 112640 =>
                  width54_xhdl57 := "011";    
                  width53_xhdl56 := "011";    
                  width52_xhdl55 := "011";    
                  width51_xhdl54 := "011";    
                  width50_xhdl53 := "011";    
                  width49_xhdl52 := "011";    
                  width48_xhdl51 := "011";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr54_xhdl333 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr53_xhdl332 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr52_xhdl331 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr51_xhdl330 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr50_xhdl329 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr49_xhdl328 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr48_xhdl327 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr53_xhdl401 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr52_xhdl400 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr51_xhdl399 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr50_xhdl398 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr49_xhdl397 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr48_xhdl396 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData54_xhdl264 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData53_xhdl263 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData52_xhdl262 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData51_xhdl261 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData50_xhdl260 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData49_xhdl259 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData48_xhdl258 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1101100" |
                          "1101101" =>
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1101010" |
                          "1101011" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1101000" |
                          "1101001" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100110" |
                          "1100111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100100" |
                          "1100101" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100010" |
                          "1100011" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1101100" |
                          "1101101" =>
                              readData_xhdl1_xhdl417 := readData54(7 
                              DOWNTO 0);    
                     WHEN "1101010" |
                          "1101011" =>
                              readData_xhdl1_xhdl417 := readData53(7 
                              DOWNTO 0);    
                     WHEN "1101000" |
                          "1101001" =>
                              readData_xhdl1_xhdl417 := readData52(7 
                              DOWNTO 0);    
                     WHEN "1100110" |
                          "1100111" =>
                              readData_xhdl1_xhdl417 := readData51(7 
                              DOWNTO 0);    
                     WHEN "1100100" |
                          "1100101" =>
                              readData_xhdl1_xhdl417 := readData50(7 
                              DOWNTO 0);    
                     WHEN "1100010" |
                          "1100011" =>
                              readData_xhdl1_xhdl417 := readData49(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" =>
                              readData_xhdl1_xhdl417 := readData48(7 
                              DOWNTO 0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 114688 =>
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 116736 =>
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 118784 =>
                  width57_xhdl60 := "011";    
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr57_xhdl336 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData57_xhdl267 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1110010" |
                          "1110011" =>
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1110010" |
                          "1110011" =>
                              readData_xhdl1_xhdl417 := readData57(7 
                              DOWNTO 0);    
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 120832 =>
                  width58_xhdl61 := "011";    
                  width57_xhdl60 := "011";    
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr58_xhdl337 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr57_xhdl336 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr57_xhdl405 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData58_xhdl268 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData57_xhdl267 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1110100" |
                          "1110101" =>
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110010" |
                          "1110011" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1110100" |
                          "1110101" =>
                              readData_xhdl1_xhdl417 := readData58(7 
                              DOWNTO 0);    
                     WHEN "1110010" |
                          "1110011" =>
                              readData_xhdl1_xhdl417 := readData57(7 
                              DOWNTO 0);    
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 122880 =>
                  width59_xhdl62 := "011";    
                  width58_xhdl61 := "011";    
                  width57_xhdl60 := "011";    
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr59_xhdl338 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr58_xhdl337 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr57_xhdl336 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr58_xhdl406 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr57_xhdl405 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData59_xhdl269 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData58_xhdl268 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData57_xhdl267 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1110110" |
                          "1110111" =>
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110100" |
                          "1110101" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110010" |
                          "1110011" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1110110" |
                          "1110111" =>
                              readData_xhdl1_xhdl417 := readData59(7 
                              DOWNTO 0);    
                     WHEN "1110100" |
                          "1110101" =>
                              readData_xhdl1_xhdl417 := readData58(7 
                              DOWNTO 0);    
                     WHEN "1110010" |
                          "1110011" =>
                              readData_xhdl1_xhdl417 := readData57(7 
                              DOWNTO 0);    
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 124928 =>
                  width60_xhdl63 := "011";    
                  width59_xhdl62 := "011";    
                  width58_xhdl61 := "011";    
                  width57_xhdl60 := "011";    
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr60_xhdl339 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr59_xhdl338 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr58_xhdl337 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr57_xhdl336 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr59_xhdl407 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr58_xhdl406 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr57_xhdl405 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData60_xhdl270 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData59_xhdl269 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData58_xhdl268 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData57_xhdl267 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1111000" |
                          "1111001" =>
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110110" |
                          "1110111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110100" |
                          "1110101" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110010" |
                          "1110011" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1111000" |
                          "1111001" =>
                              readData_xhdl1_xhdl417 := readData60(7 
                              DOWNTO 0);    
                     WHEN "1110110" |
                          "1110111" =>
                              readData_xhdl1_xhdl417 := readData59(7 
                              DOWNTO 0);    
                     WHEN "1110100" |
                          "1110101" =>
                              readData_xhdl1_xhdl417 := readData58(7 
                              DOWNTO 0);    
                     WHEN "1110010" |
                          "1110011" =>
                              readData_xhdl1_xhdl417 := readData57(7 
                              DOWNTO 0);    
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 126976 =>
                  width61_xhdl64 := "011";    
                  width60_xhdl63 := "011";    
                  width59_xhdl62 := "011";    
                  width58_xhdl61 := "011";    
                  width57_xhdl60 := "011";    
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr61_xhdl340 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr60_xhdl339 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr59_xhdl338 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr58_xhdl337 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr57_xhdl336 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr60_xhdl408 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr59_xhdl407 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr58_xhdl406 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr57_xhdl405 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData61_xhdl271 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData60_xhdl270 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData59_xhdl269 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData58_xhdl268 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData57_xhdl267 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1111010" |
                          "1111011" =>
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1111000" |
                          "1111001" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110110" |
                          "1110111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110100" |
                          "1110101" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110010" |
                          "1110011" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1111010" |
                          "1111011" =>
                              readData_xhdl1_xhdl417 := readData61(7 
                              DOWNTO 0);    
                     WHEN "1111000" |
                          "1111001" =>
                              readData_xhdl1_xhdl417 := readData60(7 
                              DOWNTO 0);    
                     WHEN "1110110" |
                          "1110111" =>
                              readData_xhdl1_xhdl417 := readData59(7 
                              DOWNTO 0);    
                     WHEN "1110100" |
                          "1110101" =>
                              readData_xhdl1_xhdl417 := readData58(7 
                              DOWNTO 0);    
                     WHEN "1110010" |
                          "1110011" =>
                              readData_xhdl1_xhdl417 := readData57(7 
                              DOWNTO 0);    
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 129024 =>
                  width62_xhdl65 := "011";    
                  width61_xhdl64 := "011";    
                  width60_xhdl63 := "011";    
                  width59_xhdl62 := "011";    
                  width58_xhdl61 := "011";    
                  width57_xhdl60 := "011";    
                  width56_xhdl59 := "011";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr62_xhdl341 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr61_xhdl340 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr60_xhdl339 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr59_xhdl338 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr58_xhdl337 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr57_xhdl336 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr56_xhdl335 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr61_xhdl409 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr60_xhdl408 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr59_xhdl407 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr58_xhdl406 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr57_xhdl405 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr56_xhdl404 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData62_xhdl272 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData61_xhdl271 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData60_xhdl270 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData59_xhdl269 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData58_xhdl268 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData57_xhdl267 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData56_xhdl266 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1111100" |
                          "1111101" =>
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1111010" |
                          "1111011" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1111000" |
                          "1111001" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110110" |
                          "1110111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110100" |
                          "1110101" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110010" |
                          "1110011" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1110000" |
                          "1110001" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1111100" |
                          "1111101" =>
                              readData_xhdl1_xhdl417 := readData62(7 
                              DOWNTO 0);    
                     WHEN "1111010" |
                          "1111011" =>
                              readData_xhdl1_xhdl417 := readData61(7 
                              DOWNTO 0);    
                     WHEN "1111000" |
                          "1111001" =>
                              readData_xhdl1_xhdl417 := readData60(7 
                              DOWNTO 0);    
                     WHEN "1110110" |
                          "1110111" =>
                              readData_xhdl1_xhdl417 := readData59(7 
                              DOWNTO 0);    
                     WHEN "1110100" |
                          "1110101" =>
                              readData_xhdl1_xhdl417 := readData58(7 
                              DOWNTO 0);    
                     WHEN "1110010" |
                          "1110011" =>
                              readData_xhdl1_xhdl417 := readData57(7 
                              DOWNTO 0);    
                     WHEN "1110000" |
                          "1110001" =>
                              readData_xhdl1_xhdl417 := readData56(7 
                              DOWNTO 0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 131072 =>
                  width63_xhdl66 := "000";    
                  width62_xhdl65 := "000";    
                  width61_xhdl64 := "000";    
                  width60_xhdl63 := "000";    
                  width59_xhdl62 := "000";    
                  width58_xhdl61 := "000";    
                  width57_xhdl60 := "000";    
                  width56_xhdl59 := "000";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr63_xhdl342 := writeAddr(13 DOWNTO 0);    
                  writeAddr62_xhdl341 := writeAddr(13 DOWNTO 0);    
                  writeAddr61_xhdl340 := writeAddr(13 DOWNTO 0);    
                  writeAddr60_xhdl339 := writeAddr(13 DOWNTO 0);    
                  writeAddr59_xhdl338 := writeAddr(13 DOWNTO 0);    
                  writeAddr58_xhdl337 := writeAddr(13 DOWNTO 0);    
                  writeAddr57_xhdl336 := writeAddr(13 DOWNTO 0);    
                  writeAddr56_xhdl335 := writeAddr(13 DOWNTO 0);    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr63_xhdl411 := readAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData63_xhdl273 := "00000000000000000" & 
                  writeData(7);    
                  writeData62_xhdl272 := "00000000000000000" & 
                  writeData(6);    
                  writeData61_xhdl271 := "00000000000000000" & 
                  writeData(5);    
                  writeData60_xhdl270 := "00000000000000000" & 
                  writeData(4);    
                  writeData59_xhdl269 := "00000000000000000" & 
                  writeData(3);    
                  writeData58_xhdl268 := "00000000000000000" & 
                  writeData(2);    
                  writeData57_xhdl267 := "00000000000000000" & 
                  writeData(1);    
                  writeData56_xhdl266 := "00000000000000000" & 
                  writeData(0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(16 DOWNTO 10) IS
                     WHEN "1110000" |
                          "1110001" |
                          "1110010" |
                          "1110011" |
                          "1110100" |
                          "1110101" |
                          "1110110" |
                          "1110111" |
                          "1111000" |
                          "1111001" |
                          "1111010" |
                          "1111011" |
                          "1111100" |
                          "1111101" |
                          "1111110" |
                          "1111111" =>
                              wen_a63_xhdl135 := '0' & wen;    
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(16 DOWNTO 10) IS
                     WHEN "1110000" |
                          "1110001" |
                          "1110010" |
                          "1110011" |
                          "1110100" |
                          "1110101" |
                          "1110110" |
                          "1110111" |
                          "1111000" |
                          "1111001" |
                          "1111010" |
                          "1111011" |
                          "1111100" |
                          "1111101" |
                          "1111110" |
                          "1111111" =>
                              readData_xhdl1_xhdl417 := readData63(0) & 
                              readData62(0) & readData61(0) & 
                              readData60(0) & readData59(0) & 
                              readData58(0) & readData57(0) & 
                              readData56(0);    
                     WHEN "1100000" |
                          "1100001" |
                          "1100010" |
                          "1100011" |
                          "1100100" |
                          "1100101" |
                          "1100110" |
                          "1100111" |
                          "1101000" |
                          "1101001" |
                          "1101010" |
                          "1101011" |
                          "1101100" |
                          "1101101" |
                          "1101110" |
                          "1101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "1010000" |
                          "1010001" |
                          "1010010" |
                          "1010011" |
                          "1010100" |
                          "1010101" |
                          "1010110" |
                          "1010111" |
                          "1011000" |
                          "1011001" |
                          "1011010" |
                          "1011011" |
                          "1011100" |
                          "1011101" |
                          "1011110" |
                          "1011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "1000000" |
                          "1000001" |
                          "1000010" |
                          "1000011" |
                          "1000100" |
                          "1000101" |
                          "1000110" |
                          "1000111" |
                          "1001000" |
                          "1001001" |
                          "1001010" |
                          "1001011" |
                          "1001100" |
                          "1001101" |
                          "1001110" |
                          "1001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "0110000" |
                          "0110001" |
                          "0110010" |
                          "0110011" |
                          "0110100" |
                          "0110101" |
                          "0110110" |
                          "0110111" |
                          "0111000" |
                          "0111001" |
                          "0111010" |
                          "0111011" |
                          "0111100" |
                          "0111101" |
                          "0111110" |
                          "0111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "0100000" |
                          "0100001" |
                          "0100010" |
                          "0100011" |
                          "0100100" |
                          "0100101" |
                          "0100110" |
                          "0100111" |
                          "0101000" |
                          "0101001" |
                          "0101010" |
                          "0101011" |
                          "0101100" |
                          "0101101" |
                          "0101110" |
                          "0101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "0010000" |
                          "0010001" |
                          "0010010" |
                          "0010011" |
                          "0010100" |
                          "0010101" |
                          "0010110" |
                          "0010111" |
                          "0011000" |
                          "0011001" |
                          "0011010" |
                          "0011011" |
                          "0011100" |
                          "0011101" |
                          "0011110" |
                          "0011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "0000000" |
                          "0000001" |
                          "0000010" |
                          "0000011" |
                          "0000100" |
                          "0000101" |
                          "0000110" |
                          "0000111" |
                          "0001000" |
                          "0001001" |
                          "0001010" |
                          "0001011" |
                          "0001100" |
                          "0001101" |
                          "0001110" |
                          "0001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 133120 =>
                  width64_xhdl67 := "011";    
                  width63_xhdl66 := "000";    
                  width62_xhdl65 := "000";    
                  width61_xhdl64 := "000";    
                  width60_xhdl63 := "000";    
                  width59_xhdl62 := "000";    
                  width58_xhdl61 := "000";    
                  width57_xhdl60 := "000";    
                  width56_xhdl59 := "000";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr64_xhdl343 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr63_xhdl342 := writeAddr(13 DOWNTO 0);    
                  writeAddr62_xhdl341 := writeAddr(13 DOWNTO 0);    
                  writeAddr61_xhdl340 := writeAddr(13 DOWNTO 0);    
                  writeAddr60_xhdl339 := writeAddr(13 DOWNTO 0);    
                  writeAddr59_xhdl338 := writeAddr(13 DOWNTO 0);    
                  writeAddr58_xhdl337 := writeAddr(13 DOWNTO 0);    
                  writeAddr57_xhdl336 := writeAddr(13 DOWNTO 0);    
                  writeAddr56_xhdl335 := writeAddr(13 DOWNTO 0);    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr64_xhdl412 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr63_xhdl411 := readAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData64_xhdl274 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData63_xhdl273 := "00000000000000000" & 
                  writeData(7);    
                  writeData62_xhdl272 := "00000000000000000" & 
                  writeData(6);    
                  writeData61_xhdl271 := "00000000000000000" & 
                  writeData(5);    
                  writeData60_xhdl270 := "00000000000000000" & 
                  writeData(4);    
                  writeData59_xhdl269 := "00000000000000000" & 
                  writeData(3);    
                  writeData58_xhdl268 := "00000000000000000" & 
                  writeData(2);    
                  writeData57_xhdl267 := "00000000000000000" & 
                  writeData(1);    
                  writeData56_xhdl266 := "00000000000000000" & 
                  writeData(0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(17 DOWNTO 10) IS
                     WHEN "10000000" |
                          "10000001" =>
                              wen_a64_xhdl136 := '0' & wen;    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & wen;    
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(17 DOWNTO 10) IS
                     WHEN "10000000" |
                          "10000001" =>
                              readData_xhdl1_xhdl417 := readData64(7 
                              DOWNTO 0);    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              readData_xhdl1_xhdl417 := readData63(0) & 
                              readData62(0) & readData61(0) & 
                              readData60(0) & readData59(0) & 
                              readData58(0) & readData57(0) & 
                              readData56(0);    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 135168 =>
                  width65_xhdl68 := "011";    
                  width64_xhdl67 := "011";    
                  width63_xhdl66 := "000";    
                  width62_xhdl65 := "000";    
                  width61_xhdl64 := "000";    
                  width60_xhdl63 := "000";    
                  width59_xhdl62 := "000";    
                  width58_xhdl61 := "000";    
                  width57_xhdl60 := "000";    
                  width56_xhdl59 := "000";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr65_xhdl344 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr64_xhdl343 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr63_xhdl342 := writeAddr(13 DOWNTO 0);    
                  writeAddr62_xhdl341 := writeAddr(13 DOWNTO 0);    
                  writeAddr61_xhdl340 := writeAddr(13 DOWNTO 0);    
                  writeAddr60_xhdl339 := writeAddr(13 DOWNTO 0);    
                  writeAddr59_xhdl338 := writeAddr(13 DOWNTO 0);    
                  writeAddr58_xhdl337 := writeAddr(13 DOWNTO 0);    
                  writeAddr57_xhdl336 := writeAddr(13 DOWNTO 0);    
                  writeAddr56_xhdl335 := writeAddr(13 DOWNTO 0);    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr65_xhdl413 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr64_xhdl412 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr63_xhdl411 := readAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData65_xhdl275 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData64_xhdl274 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData63_xhdl273 := "00000000000000000" & 
                  writeData(7);    
                  writeData62_xhdl272 := "00000000000000000" & 
                  writeData(6);    
                  writeData61_xhdl271 := "00000000000000000" & 
                  writeData(5);    
                  writeData60_xhdl270 := "00000000000000000" & 
                  writeData(4);    
                  writeData59_xhdl269 := "00000000000000000" & 
                  writeData(3);    
                  writeData58_xhdl268 := "00000000000000000" & 
                  writeData(2);    
                  writeData57_xhdl267 := "00000000000000000" & 
                  writeData(1);    
                  writeData56_xhdl266 := "00000000000000000" & 
                  writeData(0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(17 DOWNTO 10) IS
                     WHEN "10000010" |
                          "10000011" =>
                              wen_a65_xhdl137 := '0' & wen;    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000000" |
                          "10000001" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & wen;    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & wen;    
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(17 DOWNTO 10) IS
                     WHEN "10000010" |
                          "10000011" =>
                              readData_xhdl1_xhdl417 := readData65(7 
                              DOWNTO 0);    
                     WHEN "10000000" |
                          "10000001" =>
                              readData_xhdl1_xhdl417 := readData64(7 
                              DOWNTO 0);    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              readData_xhdl1_xhdl417 := readData63(0) & 
                              readData62(0) & readData61(0) & 
                              readData60(0) & readData59(0) & 
                              readData58(0) & readData57(0) & 
                              readData56(0);    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 137216 =>
                  width66_xhdl69 := "011";    
                  width65_xhdl68 := "011";    
                  width64_xhdl67 := "011";    
                  width63_xhdl66 := "000";    
                  width62_xhdl65 := "000";    
                  width61_xhdl64 := "000";    
                  width60_xhdl63 := "000";    
                  width59_xhdl62 := "000";    
                  width58_xhdl61 := "000";    
                  width57_xhdl60 := "000";    
                  width56_xhdl59 := "000";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr66_xhdl345 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr65_xhdl344 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr64_xhdl343 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr63_xhdl342 := writeAddr(13 DOWNTO 0);    
                  writeAddr62_xhdl341 := writeAddr(13 DOWNTO 0);    
                  writeAddr61_xhdl340 := writeAddr(13 DOWNTO 0);    
                  writeAddr60_xhdl339 := writeAddr(13 DOWNTO 0);    
                  writeAddr59_xhdl338 := writeAddr(13 DOWNTO 0);    
                  writeAddr58_xhdl337 := writeAddr(13 DOWNTO 0);    
                  writeAddr57_xhdl336 := writeAddr(13 DOWNTO 0);    
                  writeAddr56_xhdl335 := writeAddr(13 DOWNTO 0);    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr66_xhdl414 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr65_xhdl413 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr64_xhdl412 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr63_xhdl411 := readAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData66_xhdl276 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData65_xhdl275 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData64_xhdl274 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData63_xhdl273 := "00000000000000000" & 
                  writeData(7);    
                  writeData62_xhdl272 := "00000000000000000" & 
                  writeData(6);    
                  writeData61_xhdl271 := "00000000000000000" & 
                  writeData(5);    
                  writeData60_xhdl270 := "00000000000000000" & 
                  writeData(4);    
                  writeData59_xhdl269 := "00000000000000000" & 
                  writeData(3);    
                  writeData58_xhdl268 := "00000000000000000" & 
                  writeData(2);    
                  writeData57_xhdl267 := "00000000000000000" & 
                  writeData(1);    
                  writeData56_xhdl266 := "00000000000000000" & 
                  writeData(0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(17 DOWNTO 10) IS
                     WHEN "10000100" |
                          "10000101" =>
                              wen_a66_xhdl138 := '0' & wen;    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000010" |
                          "10000011" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & wen;    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000000" |
                          "10000001" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & wen;    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & wen;    
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(17 DOWNTO 10) IS
                     WHEN "10000100" |
                          "10000101" =>
                              readData_xhdl1_xhdl417 := readData66(7 
                              DOWNTO 0);    
                     WHEN "10000010" |
                          "10000011" =>
                              readData_xhdl1_xhdl417 := readData65(7 
                              DOWNTO 0);    
                     WHEN "10000000" |
                          "10000001" =>
                              readData_xhdl1_xhdl417 := readData64(7 
                              DOWNTO 0);    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              readData_xhdl1_xhdl417 := readData63(0) & 
                              readData62(0) & readData61(0) & 
                              readData60(0) & readData59(0) & 
                              readData58(0) & readData57(0) & 
                              readData56(0);    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[17:10])
                  
                  
         WHEN 139264 =>
                  width67_xhdl70 := "011";    
                  width66_xhdl69 := "011";    
                  width65_xhdl68 := "011";    
                  width64_xhdl67 := "011";    
                  width63_xhdl66 := "000";    
                  width62_xhdl65 := "000";    
                  width61_xhdl64 := "000";    
                  width60_xhdl63 := "000";    
                  width59_xhdl62 := "000";    
                  width58_xhdl61 := "000";    
                  width57_xhdl60 := "000";    
                  width56_xhdl59 := "000";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr67_xhdl346 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr66_xhdl345 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr65_xhdl344 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr64_xhdl343 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr63_xhdl342 := writeAddr(13 DOWNTO 0);    
                  writeAddr62_xhdl341 := writeAddr(13 DOWNTO 0);    
                  writeAddr61_xhdl340 := writeAddr(13 DOWNTO 0);    
                  writeAddr60_xhdl339 := writeAddr(13 DOWNTO 0);    
                  writeAddr59_xhdl338 := writeAddr(13 DOWNTO 0);    
                  writeAddr58_xhdl337 := writeAddr(13 DOWNTO 0);    
                  writeAddr57_xhdl336 := writeAddr(13 DOWNTO 0);    
                  writeAddr56_xhdl335 := writeAddr(13 DOWNTO 0);    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr67_xhdl415 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr66_xhdl414 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr65_xhdl413 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr64_xhdl412 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr63_xhdl411 := readAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData67_xhdl277 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData66_xhdl276 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData65_xhdl275 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData64_xhdl274 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData63_xhdl273 := "00000000000000000" & 
                  writeData(7);    
                  writeData62_xhdl272 := "00000000000000000" & 
                  writeData(6);    
                  writeData61_xhdl271 := "00000000000000000" & 
                  writeData(5);    
                  writeData60_xhdl270 := "00000000000000000" & 
                  writeData(4);    
                  writeData59_xhdl269 := "00000000000000000" & 
                  writeData(3);    
                  writeData58_xhdl268 := "00000000000000000" & 
                  writeData(2);    
                  writeData57_xhdl267 := "00000000000000000" & 
                  writeData(1);    
                  writeData56_xhdl266 := "00000000000000000" & 
                  writeData(0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(17 DOWNTO 10) IS
                     WHEN "10000110" |
                          "10000111" =>
                              wen_a67_xhdl139 := '0' & wen;    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000100" |
                          "10000101" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & wen;    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000010" |
                          "10000011" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & wen;    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000000" |
                          "10000001" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & wen;    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & wen;    
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(17 DOWNTO 10) IS
                     WHEN "10000110" |
                          "10000111" =>
                              readData_xhdl1_xhdl417 := readData67(7 
                              DOWNTO 0);    
                     WHEN "10000100" |
                          "10000101" =>
                              readData_xhdl1_xhdl417 := readData66(7 
                              DOWNTO 0);    
                     WHEN "10000010" |
                          "10000011" =>
                              readData_xhdl1_xhdl417 := readData65(7 
                              DOWNTO 0);    
                     WHEN "10000000" |
                          "10000001" =>
                              readData_xhdl1_xhdl417 := readData64(7 
                              DOWNTO 0);    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              readData_xhdl1_xhdl417 := readData63(0) & 
                              readData62(0) & readData61(0) & 
                              readData60(0) & readData59(0) & 
                              readData58(0) & readData57(0) & 
                              readData56(0);    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN 141312 =>
                  width68_xhdl71 := "011";    
                  width67_xhdl70 := "011";    
                  width66_xhdl69 := "011";    
                  width65_xhdl68 := "011";    
                  width64_xhdl67 := "011";    
                  width63_xhdl66 := "000";    
                  width62_xhdl65 := "000";    
                  width61_xhdl64 := "000";    
                  width60_xhdl63 := "000";    
                  width59_xhdl62 := "000";    
                  width58_xhdl61 := "000";    
                  width57_xhdl60 := "000";    
                  width56_xhdl59 := "000";    
                  width55_xhdl58 := "000";    
                  width54_xhdl57 := "000";    
                  width53_xhdl56 := "000";    
                  width52_xhdl55 := "000";    
                  width51_xhdl54 := "000";    
                  width50_xhdl53 := "000";    
                  width49_xhdl52 := "000";    
                  width48_xhdl51 := "000";    
                  width47_xhdl50 := "000";    
                  width46_xhdl49 := "000";    
                  width45_xhdl48 := "000";    
                  width44_xhdl47 := "000";    
                  width43_xhdl46 := "000";    
                  width42_xhdl45 := "000";    
                  width41_xhdl44 := "000";    
                  width40_xhdl43 := "000";    
                  width39_xhdl42 := "000";    
                  width38_xhdl41 := "000";    
                  width37_xhdl40 := "000";    
                  width36_xhdl39 := "000";    
                  width35_xhdl38 := "000";    
                  width34_xhdl37 := "000";    
                  width33_xhdl36 := "000";    
                  width32_xhdl35 := "000";    
                  width31_xhdl34 := "000";    
                  width30_xhdl33 := "000";    
                  width29_xhdl32 := "000";    
                  width28_xhdl31 := "000";    
                  width27_xhdl30 := "000";    
                  width26_xhdl29 := "000";    
                  width25_xhdl28 := "000";    
                  width24_xhdl27 := "000";    
                  width23_xhdl26 := "000";    
                  width22_xhdl25 := "000";    
                  width21_xhdl24 := "000";    
                  width20_xhdl23 := "000";    
                  width19_xhdl22 := "000";    
                  width18_xhdl21 := "000";    
                  width17_xhdl20 := "000";    
                  width16_xhdl19 := "000";    
                  width15_xhdl18 := "000";    
                  width14_xhdl17 := "000";    
                  width13_xhdl16 := "000";    
                  width12_xhdl15 := "000";    
                  width11_xhdl14 := "000";    
                  width10_xhdl13 := "000";    
                  width9_xhdl12 := "000";    
                  width8_xhdl11 := "000";    
                  width7_xhdl10 := "000";    
                  width6_xhdl9 := "000";    
                  width5_xhdl8 := "000";    
                  width4_xhdl7 := "000";    
                  width3_xhdl6 := "000";    
                  width2_xhdl5 := "000";    
                  width1_xhdl4 := "000";    
                  width0_xhdl3 := "000";    
                  writeAddr68_xhdl347 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr67_xhdl346 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr66_xhdl345 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr65_xhdl344 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr64_xhdl343 := writeAddr(10 DOWNTO 0) & "000"; 
                  writeAddr63_xhdl342 := writeAddr(13 DOWNTO 0);    
                  writeAddr62_xhdl341 := writeAddr(13 DOWNTO 0);    
                  writeAddr61_xhdl340 := writeAddr(13 DOWNTO 0);    
                  writeAddr60_xhdl339 := writeAddr(13 DOWNTO 0);    
                  writeAddr59_xhdl338 := writeAddr(13 DOWNTO 0);    
                  writeAddr58_xhdl337 := writeAddr(13 DOWNTO 0);    
                  writeAddr57_xhdl336 := writeAddr(13 DOWNTO 0);    
                  writeAddr56_xhdl335 := writeAddr(13 DOWNTO 0);    
                  writeAddr55_xhdl334 := writeAddr(13 DOWNTO 0);    
                  writeAddr54_xhdl333 := writeAddr(13 DOWNTO 0);    
                  writeAddr53_xhdl332 := writeAddr(13 DOWNTO 0);    
                  writeAddr52_xhdl331 := writeAddr(13 DOWNTO 0);    
                  writeAddr51_xhdl330 := writeAddr(13 DOWNTO 0);    
                  writeAddr50_xhdl329 := writeAddr(13 DOWNTO 0);    
                  writeAddr49_xhdl328 := writeAddr(13 DOWNTO 0);    
                  writeAddr48_xhdl327 := writeAddr(13 DOWNTO 0);    
                  writeAddr47_xhdl326 := writeAddr(13 DOWNTO 0);    
                  writeAddr46_xhdl325 := writeAddr(13 DOWNTO 0);    
                  writeAddr45_xhdl324 := writeAddr(13 DOWNTO 0);    
                  writeAddr44_xhdl323 := writeAddr(13 DOWNTO 0);    
                  writeAddr43_xhdl322 := writeAddr(13 DOWNTO 0);    
                  writeAddr42_xhdl321 := writeAddr(13 DOWNTO 0);    
                  writeAddr41_xhdl320 := writeAddr(13 DOWNTO 0);    
                  writeAddr40_xhdl319 := writeAddr(13 DOWNTO 0);    
                  writeAddr39_xhdl318 := writeAddr(13 DOWNTO 0);    
                  writeAddr38_xhdl317 := writeAddr(13 DOWNTO 0);    
                  writeAddr37_xhdl316 := writeAddr(13 DOWNTO 0);    
                  writeAddr36_xhdl315 := writeAddr(13 DOWNTO 0);    
                  writeAddr35_xhdl314 := writeAddr(13 DOWNTO 0);    
                  writeAddr34_xhdl313 := writeAddr(13 DOWNTO 0);    
                  writeAddr33_xhdl312 := writeAddr(13 DOWNTO 0);    
                  writeAddr32_xhdl311 := writeAddr(13 DOWNTO 0);    
                  writeAddr31_xhdl310 := writeAddr(13 DOWNTO 0);    
                  writeAddr30_xhdl309 := writeAddr(13 DOWNTO 0);    
                  writeAddr29_xhdl308 := writeAddr(13 DOWNTO 0);    
                  writeAddr28_xhdl307 := writeAddr(13 DOWNTO 0);    
                  writeAddr27_xhdl306 := writeAddr(13 DOWNTO 0);    
                  writeAddr26_xhdl305 := writeAddr(13 DOWNTO 0);    
                  writeAddr25_xhdl304 := writeAddr(13 DOWNTO 0);    
                  writeAddr24_xhdl303 := writeAddr(13 DOWNTO 0);    
                  writeAddr23_xhdl302 := writeAddr(13 DOWNTO 0);    
                  writeAddr22_xhdl301 := writeAddr(13 DOWNTO 0);    
                  writeAddr21_xhdl300 := writeAddr(13 DOWNTO 0);    
                  writeAddr20_xhdl299 := writeAddr(13 DOWNTO 0);    
                  writeAddr19_xhdl298 := writeAddr(13 DOWNTO 0);    
                  writeAddr18_xhdl297 := writeAddr(13 DOWNTO 0);    
                  writeAddr17_xhdl296 := writeAddr(13 DOWNTO 0);    
                  writeAddr16_xhdl295 := writeAddr(13 DOWNTO 0);    
                  writeAddr15_xhdl294 := writeAddr(13 DOWNTO 0);    
                  writeAddr14_xhdl293 := writeAddr(13 DOWNTO 0);    
                  writeAddr13_xhdl292 := writeAddr(13 DOWNTO 0);    
                  writeAddr12_xhdl291 := writeAddr(13 DOWNTO 0);    
                  writeAddr11_xhdl290 := writeAddr(13 DOWNTO 0);    
                  writeAddr10_xhdl289 := writeAddr(13 DOWNTO 0);    
                  writeAddr9_xhdl288 := writeAddr(13 DOWNTO 0);    
                  writeAddr8_xhdl287 := writeAddr(13 DOWNTO 0);    
                  writeAddr7_xhdl286 := writeAddr(13 DOWNTO 0);    
                  writeAddr6_xhdl285 := writeAddr(13 DOWNTO 0);    
                  writeAddr5_xhdl284 := writeAddr(13 DOWNTO 0);    
                  writeAddr4_xhdl283 := writeAddr(13 DOWNTO 0);    
                  writeAddr3_xhdl282 := writeAddr(13 DOWNTO 0);    
                  writeAddr2_xhdl281 := writeAddr(13 DOWNTO 0);    
                  writeAddr1_xhdl280 := writeAddr(13 DOWNTO 0);    
                  writeAddr0_xhdl279 := writeAddr(13 DOWNTO 0);    
                  readAddr68_xhdl416 := readAddr(10 DOWNTO 0) & "000"; 
                  readAddr67_xhdl415 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr66_xhdl414 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr65_xhdl413 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr64_xhdl412 := readAddr(10 DOWNTO 0) & "000";   
                  readAddr63_xhdl411 := readAddr(13 DOWNTO 0);    
                  readAddr62_xhdl410 := readAddr(13 DOWNTO 0);    
                  readAddr61_xhdl409 := readAddr(13 DOWNTO 0);    
                  readAddr60_xhdl408 := readAddr(13 DOWNTO 0);    
                  readAddr59_xhdl407 := readAddr(13 DOWNTO 0);    
                  readAddr58_xhdl406 := readAddr(13 DOWNTO 0);    
                  readAddr57_xhdl405 := readAddr(13 DOWNTO 0);    
                  readAddr56_xhdl404 := readAddr(13 DOWNTO 0);    
                  readAddr55_xhdl403 := readAddr(13 DOWNTO 0);    
                  readAddr54_xhdl402 := readAddr(13 DOWNTO 0);    
                  readAddr53_xhdl401 := readAddr(13 DOWNTO 0);    
                  readAddr52_xhdl400 := readAddr(13 DOWNTO 0);    
                  readAddr51_xhdl399 := readAddr(13 DOWNTO 0);    
                  readAddr50_xhdl398 := readAddr(13 DOWNTO 0);    
                  readAddr49_xhdl397 := readAddr(13 DOWNTO 0);    
                  readAddr48_xhdl396 := readAddr(13 DOWNTO 0);    
                  readAddr47_xhdl395 := readAddr(13 DOWNTO 0);    
                  readAddr46_xhdl394 := readAddr(13 DOWNTO 0);    
                  readAddr45_xhdl393 := readAddr(13 DOWNTO 0);    
                  readAddr44_xhdl392 := readAddr(13 DOWNTO 0);    
                  readAddr43_xhdl391 := readAddr(13 DOWNTO 0);    
                  readAddr42_xhdl390 := readAddr(13 DOWNTO 0);    
                  readAddr41_xhdl389 := readAddr(13 DOWNTO 0);    
                  readAddr40_xhdl388 := readAddr(13 DOWNTO 0);    
                  readAddr39_xhdl387 := readAddr(13 DOWNTO 0);    
                  readAddr38_xhdl386 := readAddr(13 DOWNTO 0);    
                  readAddr37_xhdl385 := readAddr(13 DOWNTO 0);    
                  readAddr36_xhdl384 := readAddr(13 DOWNTO 0);    
                  readAddr35_xhdl383 := readAddr(13 DOWNTO 0);    
                  readAddr34_xhdl382 := readAddr(13 DOWNTO 0);    
                  readAddr33_xhdl381 := readAddr(13 DOWNTO 0);    
                  readAddr32_xhdl380 := readAddr(13 DOWNTO 0);    
                  readAddr31_xhdl379 := readAddr(13 DOWNTO 0);    
                  readAddr30_xhdl378 := readAddr(13 DOWNTO 0);    
                  readAddr29_xhdl377 := readAddr(13 DOWNTO 0);    
                  readAddr28_xhdl376 := readAddr(13 DOWNTO 0);    
                  readAddr27_xhdl375 := readAddr(13 DOWNTO 0);    
                  readAddr26_xhdl374 := readAddr(13 DOWNTO 0);    
                  readAddr25_xhdl373 := readAddr(13 DOWNTO 0);    
                  readAddr24_xhdl372 := readAddr(13 DOWNTO 0);    
                  readAddr23_xhdl371 := readAddr(13 DOWNTO 0);    
                  readAddr22_xhdl370 := readAddr(13 DOWNTO 0);    
                  readAddr21_xhdl369 := readAddr(13 DOWNTO 0);    
                  readAddr20_xhdl368 := readAddr(13 DOWNTO 0);    
                  readAddr19_xhdl367 := readAddr(13 DOWNTO 0);    
                  readAddr18_xhdl366 := readAddr(13 DOWNTO 0);    
                  readAddr17_xhdl365 := readAddr(13 DOWNTO 0);    
                  readAddr16_xhdl364 := readAddr(13 DOWNTO 0);    
                  readAddr15_xhdl363 := readAddr(13 DOWNTO 0);    
                  readAddr14_xhdl362 := readAddr(13 DOWNTO 0);    
                  readAddr13_xhdl361 := readAddr(13 DOWNTO 0);    
                  readAddr12_xhdl360 := readAddr(13 DOWNTO 0);    
                  readAddr11_xhdl359 := readAddr(13 DOWNTO 0);    
                  readAddr10_xhdl358 := readAddr(13 DOWNTO 0);    
                  readAddr9_xhdl357 := readAddr(13 DOWNTO 0);    
                  readAddr8_xhdl356 := readAddr(13 DOWNTO 0);    
                  readAddr7_xhdl355 := readAddr(13 DOWNTO 0);    
                  readAddr6_xhdl354 := readAddr(13 DOWNTO 0);    
                  readAddr5_xhdl353 := readAddr(13 DOWNTO 0);    
                  readAddr4_xhdl352 := readAddr(13 DOWNTO 0);    
                  readAddr3_xhdl351 := readAddr(13 DOWNTO 0);    
                  readAddr2_xhdl350 := readAddr(13 DOWNTO 0);    
                  readAddr1_xhdl349 := readAddr(13 DOWNTO 0);    
                  readAddr0_xhdl348 := readAddr(13 DOWNTO 0);    
                  writeData68_xhdl278 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData67_xhdl277 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData66_xhdl276 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData65_xhdl275 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData64_xhdl274 := "0000000000" & writeData(7 
                  DOWNTO 0);    
                  writeData63_xhdl273 := "00000000000000000" & 
                  writeData(7);    
                  writeData62_xhdl272 := "00000000000000000" & 
                  writeData(6);    
                  writeData61_xhdl271 := "00000000000000000" & 
                  writeData(5);    
                  writeData60_xhdl270 := "00000000000000000" & 
                  writeData(4);    
                  writeData59_xhdl269 := "00000000000000000" & 
                  writeData(3);    
                  writeData58_xhdl268 := "00000000000000000" & 
                  writeData(2);    
                  writeData57_xhdl267 := "00000000000000000" & 
                  writeData(1);    
                  writeData56_xhdl266 := "00000000000000000" & 
                  writeData(0);    
                  writeData55_xhdl265 := "00000000000000000" & 
                  writeData(7);    
                  writeData54_xhdl264 := "00000000000000000" & 
                  writeData(6);    
                  writeData53_xhdl263 := "00000000000000000" & 
                  writeData(5);    
                  writeData52_xhdl262 := "00000000000000000" & 
                  writeData(4);    
                  writeData51_xhdl261 := "00000000000000000" & 
                  writeData(3);    
                  writeData50_xhdl260 := "00000000000000000" & 
                  writeData(2);    
                  writeData49_xhdl259 := "00000000000000000" & 
                  writeData(1);    
                  writeData48_xhdl258 := "00000000000000000" & 
                  writeData(0);    
                  writeData47_xhdl257 := "00000000000000000" & 
                  writeData(7);    
                  writeData46_xhdl256 := "00000000000000000" & 
                  writeData(6);    
                  writeData45_xhdl255 := "00000000000000000" & 
                  writeData(5);    
                  writeData44_xhdl254 := "00000000000000000" & 
                  writeData(4);    
                  writeData43_xhdl253 := "00000000000000000" & 
                  writeData(3);    
                  writeData42_xhdl252 := "00000000000000000" & 
                  writeData(2);    
                  writeData41_xhdl251 := "00000000000000000" & 
                  writeData(1);    
                  writeData40_xhdl250 := "00000000000000000" & 
                  writeData(0);    
                  writeData39_xhdl249 := "00000000000000000" & 
                  writeData(7);    
                  writeData38_xhdl248 := "00000000000000000" & 
                  writeData(6);    
                  writeData37_xhdl247 := "00000000000000000" & 
                  writeData(5);    
                  writeData36_xhdl246 := "00000000000000000" & 
                  writeData(4);    
                  writeData35_xhdl245 := "00000000000000000" & 
                  writeData(3);    
                  writeData34_xhdl244 := "00000000000000000" & 
                  writeData(2);    
                  writeData33_xhdl243 := "00000000000000000" & 
                  writeData(1);    
                  writeData32_xhdl242 := "00000000000000000" & 
                  writeData(0);    
                  writeData31_xhdl241 := "00000000000000000" & 
                  writeData(7);    
                  writeData30_xhdl240 := "00000000000000000" & 
                  writeData(6);    
                  writeData29_xhdl239 := "00000000000000000" & 
                  writeData(5);    
                  writeData28_xhdl238 := "00000000000000000" & 
                  writeData(4);    
                  writeData27_xhdl237 := "00000000000000000" & 
                  writeData(3);    
                  writeData26_xhdl236 := "00000000000000000" & 
                  writeData(2);    
                  writeData25_xhdl235 := "00000000000000000" & 
                  writeData(1);    
                  writeData24_xhdl234 := "00000000000000000" & 
                  writeData(0);    
                  writeData23_xhdl233 := "00000000000000000" & 
                  writeData(7);    
                  writeData22_xhdl232 := "00000000000000000" & 
                  writeData(6);    
                  writeData21_xhdl231 := "00000000000000000" & 
                  writeData(5);    
                  writeData20_xhdl230 := "00000000000000000" & 
                  writeData(4);    
                  writeData19_xhdl229 := "00000000000000000" & 
                  writeData(3);    
                  writeData18_xhdl228 := "00000000000000000" & 
                  writeData(2);    
                  writeData17_xhdl227 := "00000000000000000" & 
                  writeData(1);    
                  writeData16_xhdl226 := "00000000000000000" & 
                  writeData(0);    
                  writeData15_xhdl225 := "00000000000000000" & 
                  writeData(7);    
                  writeData14_xhdl224 := "00000000000000000" & 
                  writeData(6);    
                  writeData13_xhdl223 := "00000000000000000" & 
                  writeData(5);    
                  writeData12_xhdl222 := "00000000000000000" & 
                  writeData(4);    
                  writeData11_xhdl221 := "00000000000000000" & 
                  writeData(3);    
                  writeData10_xhdl220 := "00000000000000000" & 
                  writeData(2);    
                  writeData9_xhdl219 := "00000000000000000" & 
                  writeData(1);    
                  writeData8_xhdl218 := "00000000000000000" & 
                  writeData(0);    
                  writeData7_xhdl217 := "00000000000000000" & 
                  writeData(7);    
                  writeData6_xhdl216 := "00000000000000000" & 
                  writeData(6);    
                  writeData5_xhdl215 := "00000000000000000" & 
                  writeData(5);    
                  writeData4_xhdl214 := "00000000000000000" & 
                  writeData(4);    
                  writeData3_xhdl213 := "00000000000000000" & 
                  writeData(3);    
                  writeData2_xhdl212 := "00000000000000000" & 
                  writeData(2);    
                  writeData1_xhdl211 := "00000000000000000" & 
                  writeData(1);    
                  writeData0_xhdl210 := "00000000000000000" & 
                  writeData(0);    
                  CASE writeAddr(17 DOWNTO 10) IS
                     WHEN "10001000" |
                          "10001001" =>
                              wen_a68_xhdl140 := '0' & wen;    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000110" |
                          "10000111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & wen;    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000100" |
                          "10000101" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & wen;    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000010" |
                          "10000011" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & wen;    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "10000000" |
                          "10000001" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & wen;    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & wen;    
                              wen_a62_xhdl134 := '0' & wen;    
                              wen_a61_xhdl133 := '0' & wen;    
                              wen_a60_xhdl132 := '0' & wen;    
                              wen_a59_xhdl131 := '0' & wen;    
                              wen_a58_xhdl130 := '0' & wen;    
                              wen_a57_xhdl129 := '0' & wen;    
                              wen_a56_xhdl128 := '0' & wen;    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & wen;    
                              wen_a54_xhdl126 := '0' & wen;    
                              wen_a53_xhdl125 := '0' & wen;    
                              wen_a52_xhdl124 := '0' & wen;    
                              wen_a51_xhdl123 := '0' & wen;    
                              wen_a50_xhdl122 := '0' & wen;    
                              wen_a49_xhdl121 := '0' & wen;    
                              wen_a48_xhdl120 := '0' & wen;    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & wen;    
                              wen_a46_xhdl118 := '0' & wen;    
                              wen_a45_xhdl117 := '0' & wen;    
                              wen_a44_xhdl116 := '0' & wen;    
                              wen_a43_xhdl115 := '0' & wen;    
                              wen_a42_xhdl114 := '0' & wen;    
                              wen_a41_xhdl113 := '0' & wen;    
                              wen_a40_xhdl112 := '0' & wen;    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & wen;    
                              wen_a38_xhdl110 := '0' & wen;    
                              wen_a37_xhdl109 := '0' & wen;    
                              wen_a36_xhdl108 := '0' & wen;    
                              wen_a35_xhdl107 := '0' & wen;    
                              wen_a34_xhdl106 := '0' & wen;    
                              wen_a33_xhdl105 := '0' & wen;    
                              wen_a32_xhdl104 := '0' & wen;    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & wen;    
                              wen_a30_xhdl102 := '0' & wen;    
                              wen_a29_xhdl101 := '0' & wen;    
                              wen_a28_xhdl100 := '0' & wen;    
                              wen_a27_xhdl99 := '0' & wen;    
                              wen_a26_xhdl98 := '0' & wen;    
                              wen_a25_xhdl97 := '0' & wen;    
                              wen_a24_xhdl96 := '0' & wen;    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & wen;    
                              wen_a22_xhdl94 := '0' & wen;    
                              wen_a21_xhdl93 := '0' & wen;    
                              wen_a20_xhdl92 := '0' & wen;    
                              wen_a19_xhdl91 := '0' & wen;    
                              wen_a18_xhdl90 := '0' & wen;    
                              wen_a17_xhdl89 := '0' & wen;    
                              wen_a16_xhdl88 := '0' & wen;    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & wen;    
                              wen_a14_xhdl86 := '0' & wen;    
                              wen_a13_xhdl85 := '0' & wen;    
                              wen_a12_xhdl84 := '0' & wen;    
                              wen_a11_xhdl83 := '0' & wen;    
                              wen_a10_xhdl82 := '0' & wen;    
                              wen_a9_xhdl81 := '0' & wen;    
                              wen_a8_xhdl80 := '0' & wen;    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & wen;    
                              wen_a6_xhdl78 := '0' & wen;    
                              wen_a5_xhdl77 := '0' & wen;    
                              wen_a4_xhdl76 := '0' & wen;    
                              wen_a3_xhdl75 := '0' & wen;    
                              wen_a2_xhdl74 := '0' & wen;    
                              wen_a1_xhdl73 := '0' & wen;    
                              wen_a0_xhdl72 := '0' & wen;    
                     WHEN OTHERS  =>
                              wen_a68_xhdl140 := '0' & '0';    
                              wen_a67_xhdl139 := '0' & '0';    
                              wen_a66_xhdl138 := '0' & '0';    
                              wen_a65_xhdl137 := '0' & '0';    
                              wen_a64_xhdl136 := '0' & '0';    
                              wen_a63_xhdl135 := '0' & '0';    
                              wen_a62_xhdl134 := '0' & '0';    
                              wen_a61_xhdl133 := '0' & '0';    
                              wen_a60_xhdl132 := '0' & '0';    
                              wen_a59_xhdl131 := '0' & '0';    
                              wen_a58_xhdl130 := '0' & '0';    
                              wen_a57_xhdl129 := '0' & '0';    
                              wen_a56_xhdl128 := '0' & '0';    
                              wen_a55_xhdl127 := '0' & '0';    
                              wen_a54_xhdl126 := '0' & '0';    
                              wen_a53_xhdl125 := '0' & '0';    
                              wen_a52_xhdl124 := '0' & '0';    
                              wen_a51_xhdl123 := '0' & '0';    
                              wen_a50_xhdl122 := '0' & '0';    
                              wen_a49_xhdl121 := '0' & '0';    
                              wen_a48_xhdl120 := '0' & '0';    
                              wen_a47_xhdl119 := '0' & '0';    
                              wen_a46_xhdl118 := '0' & '0';    
                              wen_a45_xhdl117 := '0' & '0';    
                              wen_a44_xhdl116 := '0' & '0';    
                              wen_a43_xhdl115 := '0' & '0';    
                              wen_a42_xhdl114 := '0' & '0';    
                              wen_a41_xhdl113 := '0' & '0';    
                              wen_a40_xhdl112 := '0' & '0';    
                              wen_a39_xhdl111 := '0' & '0';    
                              wen_a38_xhdl110 := '0' & '0';    
                              wen_a37_xhdl109 := '0' & '0';    
                              wen_a36_xhdl108 := '0' & '0';    
                              wen_a35_xhdl107 := '0' & '0';    
                              wen_a34_xhdl106 := '0' & '0';    
                              wen_a33_xhdl105 := '0' & '0';    
                              wen_a32_xhdl104 := '0' & '0';    
                              wen_a31_xhdl103 := '0' & '0';    
                              wen_a30_xhdl102 := '0' & '0';    
                              wen_a29_xhdl101 := '0' & '0';    
                              wen_a28_xhdl100 := '0' & '0';    
                              wen_a27_xhdl99 := '0' & '0';    
                              wen_a26_xhdl98 := '0' & '0';    
                              wen_a25_xhdl97 := '0' & '0';    
                              wen_a24_xhdl96 := '0' & '0';    
                              wen_a23_xhdl95 := '0' & '0';    
                              wen_a22_xhdl94 := '0' & '0';    
                              wen_a21_xhdl93 := '0' & '0';    
                              wen_a20_xhdl92 := '0' & '0';    
                              wen_a19_xhdl91 := '0' & '0';    
                              wen_a18_xhdl90 := '0' & '0';    
                              wen_a17_xhdl89 := '0' & '0';    
                              wen_a16_xhdl88 := '0' & '0';    
                              wen_a15_xhdl87 := '0' & '0';    
                              wen_a14_xhdl86 := '0' & '0';    
                              wen_a13_xhdl85 := '0' & '0';    
                              wen_a12_xhdl84 := '0' & '0';    
                              wen_a11_xhdl83 := '0' & '0';    
                              wen_a10_xhdl82 := '0' & '0';    
                              wen_a9_xhdl81 := '0' & '0';    
                              wen_a8_xhdl80 := '0' & '0';    
                              wen_a7_xhdl79 := '0' & '0';    
                              wen_a6_xhdl78 := '0' & '0';    
                              wen_a5_xhdl77 := '0' & '0';    
                              wen_a4_xhdl76 := '0' & '0';    
                              wen_a3_xhdl75 := '0' & '0';    
                              wen_a2_xhdl74 := '0' & '0';    
                              wen_a1_xhdl73 := '0' & '0';    
                              wen_a0_xhdl72 := '0' & '0';    
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  CASE ckRdAddr(17 DOWNTO 10) IS
                     WHEN "10001000" |
                          "10001001" =>
                              readData_xhdl1_xhdl417 := readData68(7 
                              DOWNTO 0);    
                     WHEN "10000110" |
                          "10000111" =>
                              readData_xhdl1_xhdl417 := readData67(7 
                              DOWNTO 0);    
                     WHEN "10000100" |
                          "10000101" =>
                              readData_xhdl1_xhdl417 := readData66(7 
                              DOWNTO 0);    
                     WHEN "10000010" |
                          "10000011" =>
                              readData_xhdl1_xhdl417 := readData65(7 
                              DOWNTO 0);    
                     WHEN "10000000" |
                          "10000001" =>
                              readData_xhdl1_xhdl417 := readData64(7 
                              DOWNTO 0);    
                     WHEN "01110000" |
                          "01110001" |
                          "01110010" |
                          "01110011" |
                          "01110100" |
                          "01110101" |
                          "01110110" |
                          "01110111" |
                          "01111000" |
                          "01111001" |
                          "01111010" |
                          "01111011" |
                          "01111100" |
                          "01111101" |
                          "01111110" |
                          "01111111" =>
                              readData_xhdl1_xhdl417 := readData63(0) & 
                              readData62(0) & readData61(0) & 
                              readData60(0) & readData59(0) & 
                              readData58(0) & readData57(0) & 
                              readData56(0);    
                     WHEN "01100000" |
                          "01100001" |
                          "01100010" |
                          "01100011" |
                          "01100100" |
                          "01100101" |
                          "01100110" |
                          "01100111" |
                          "01101000" |
                          "01101001" |
                          "01101010" |
                          "01101011" |
                          "01101100" |
                          "01101101" |
                          "01101110" |
                          "01101111" =>
                              readData_xhdl1_xhdl417 := readData55(0) & 
                              readData54(0) & readData53(0) & 
                              readData52(0) & readData51(0) & 
                              readData50(0) & readData49(0) & 
                              readData48(0);    
                     WHEN "01010000" |
                          "01010001" |
                          "01010010" |
                          "01010011" |
                          "01010100" |
                          "01010101" |
                          "01010110" |
                          "01010111" |
                          "01011000" |
                          "01011001" |
                          "01011010" |
                          "01011011" |
                          "01011100" |
                          "01011101" |
                          "01011110" |
                          "01011111" =>
                              readData_xhdl1_xhdl417 := readData47(0) & 
                              readData46(0) & readData45(0) & 
                              readData44(0) & readData43(0) & 
                              readData42(0) & readData41(0) & 
                              readData40(0);    
                     WHEN "01000000" |
                          "01000001" |
                          "01000010" |
                          "01000011" |
                          "01000100" |
                          "01000101" |
                          "01000110" |
                          "01000111" |
                          "01001000" |
                          "01001001" |
                          "01001010" |
                          "01001011" |
                          "01001100" |
                          "01001101" |
                          "01001110" |
                          "01001111" =>
                              readData_xhdl1_xhdl417 := readData39(0) & 
                              readData38(0) & readData37(0) & 
                              readData36(0) & readData35(0) & 
                              readData34(0) & readData33(0) & 
                              readData32(0);    
                     WHEN "00110000" |
                          "00110001" |
                          "00110010" |
                          "00110011" |
                          "00110100" |
                          "00110101" |
                          "00110110" |
                          "00110111" |
                          "00111000" |
                          "00111001" |
                          "00111010" |
                          "00111011" |
                          "00111100" |
                          "00111101" |
                          "00111110" |
                          "00111111" =>
                              readData_xhdl1_xhdl417 := readData31(0) & 
                              readData30(0) & readData29(0) & 
                              readData28(0) & readData27(0) & 
                              readData26(0) & readData25(0) & 
                              readData24(0);    
                     WHEN "00100000" |
                          "00100001" |
                          "00100010" |
                          "00100011" |
                          "00100100" |
                          "00100101" |
                          "00100110" |
                          "00100111" |
                          "00101000" |
                          "00101001" |
                          "00101010" |
                          "00101011" |
                          "00101100" |
                          "00101101" |
                          "00101110" |
                          "00101111" =>
                              readData_xhdl1_xhdl417 := readData23(0) & 
                              readData22(0) & readData21(0) & 
                              readData20(0) & readData19(0) & 
                              readData18(0) & readData17(0) & 
                              readData16(0);    
                     WHEN "00010000" |
                          "00010001" |
                          "00010010" |
                          "00010011" |
                          "00010100" |
                          "00010101" |
                          "00010110" |
                          "00010111" |
                          "00011000" |
                          "00011001" |
                          "00011010" |
                          "00011011" |
                          "00011100" |
                          "00011101" |
                          "00011110" |
                          "00011111" =>
                              readData_xhdl1_xhdl417 := readData15(0) & 
                              readData14(0) & readData13(0) & 
                              readData12(0) & readData11(0) & 
                              readData10(0) & readData9(0) & readData8(0)
                              ;    
                     WHEN "00000000" |
                          "00000001" |
                          "00000010" |
                          "00000011" |
                          "00000100" |
                          "00000101" |
                          "00000110" |
                          "00000111" |
                          "00001000" |
                          "00001001" |
                          "00001010" |
                          "00001011" |
                          "00001100" |
                          "00001101" |
                          "00001110" |
                          "00001111" =>
                              readData_xhdl1_xhdl417 := readData7(0) & 
                              readData6(0) & readData5(0) & readData4(0) 
                              & readData3(0) & readData2(0) & 
                              readData1(0) & readData0(0);    
                     WHEN OTHERS  =>
                              readData_xhdl1_xhdl417 := (OTHERS => '0'); 
                     
                  END CASE;
                  -- case (writeAddr[16:10])
                  
                  
         WHEN OTHERS =>
                  NULL;
         
         -- case: 141312
         
      END CASE;
      -- case (DEPTH)
      
      
      width0 <= width0_xhdl3;
      width1 <= width1_xhdl4;
      width2 <= width2_xhdl5;
      width3 <= width3_xhdl6;
      width4 <= width4_xhdl7;
      width5 <= width5_xhdl8;
      width6 <= width6_xhdl9;
      width7 <= width7_xhdl10;
      width8 <= width8_xhdl11;
      width9 <= width9_xhdl12;
      width10 <= width10_xhdl13;
      width11 <= width11_xhdl14;
      width12 <= width12_xhdl15;
      width13 <= width13_xhdl16;
      width14 <= width14_xhdl17;
      width15 <= width15_xhdl18;
      width16 <= width16_xhdl19;
      width17 <= width17_xhdl20;
      width18 <= width18_xhdl21;
      width19 <= width19_xhdl22;
      width20 <= width20_xhdl23;
      width21 <= width21_xhdl24;
      width22 <= width22_xhdl25;
      width23 <= width23_xhdl26;
      width24 <= width24_xhdl27;
      width25 <= width25_xhdl28;
      width26 <= width26_xhdl29;
      width27 <= width27_xhdl30;
      width28 <= width28_xhdl31;
      width29 <= width29_xhdl32;
      width30 <= width30_xhdl33;
      width31 <= width31_xhdl34;
      width32 <= width32_xhdl35;
      width33 <= width33_xhdl36;
      width34 <= width34_xhdl37;
      width35 <= width35_xhdl38;
      width36 <= width36_xhdl39;
      width37 <= width37_xhdl40;
      width38 <= width38_xhdl41;
      width39 <= width39_xhdl42;
      width40 <= width40_xhdl43;
      width41 <= width41_xhdl44;
      width42 <= width42_xhdl45;
      width43 <= width43_xhdl46;
      width44 <= width44_xhdl47;
      width45 <= width45_xhdl48;
      width46 <= width46_xhdl49;
      width47 <= width47_xhdl50;
      width48 <= width48_xhdl51;
      width49 <= width49_xhdl52;
      width50 <= width50_xhdl53;
      width51 <= width51_xhdl54;
      width52 <= width52_xhdl55;
      width53 <= width53_xhdl56;
      width54 <= width54_xhdl57;
      width55 <= width55_xhdl58;
      width56 <= width56_xhdl59;
      width57 <= width57_xhdl60;
      width58 <= width58_xhdl61;
      width59 <= width59_xhdl62;
      width60 <= width60_xhdl63;
      width61 <= width61_xhdl64;
      width62 <= width62_xhdl65;
      width63 <= width63_xhdl66;
      width64 <= width64_xhdl67;
      width65 <= width65_xhdl68;
      width66 <= width66_xhdl69;
      width67 <= width67_xhdl70;
      width68 <= width68_xhdl71;
      wen_a0 <= wen_a0_xhdl72;
      wen_a1 <= wen_a1_xhdl73;
      wen_a2 <= wen_a2_xhdl74;
      wen_a3 <= wen_a3_xhdl75;
      wen_a4 <= wen_a4_xhdl76;
      wen_a5 <= wen_a5_xhdl77;
      wen_a6 <= wen_a6_xhdl78;
      wen_a7 <= wen_a7_xhdl79;
      wen_a8 <= wen_a8_xhdl80;
      wen_a9 <= wen_a9_xhdl81;
      wen_a10 <= wen_a10_xhdl82;
      wen_a11 <= wen_a11_xhdl83;
      wen_a12 <= wen_a12_xhdl84;
      wen_a13 <= wen_a13_xhdl85;
      wen_a14 <= wen_a14_xhdl86;
      wen_a15 <= wen_a15_xhdl87;
      wen_a16 <= wen_a16_xhdl88;
      wen_a17 <= wen_a17_xhdl89;
      wen_a18 <= wen_a18_xhdl90;
      wen_a19 <= wen_a19_xhdl91;
      wen_a20 <= wen_a20_xhdl92;
      wen_a21 <= wen_a21_xhdl93;
      wen_a22 <= wen_a22_xhdl94;
      wen_a23 <= wen_a23_xhdl95;
      wen_a24 <= wen_a24_xhdl96;
      wen_a25 <= wen_a25_xhdl97;
      wen_a26 <= wen_a26_xhdl98;
      wen_a27 <= wen_a27_xhdl99;
      wen_a28 <= wen_a28_xhdl100;
      wen_a29 <= wen_a29_xhdl101;
      wen_a30 <= wen_a30_xhdl102;
      wen_a31 <= wen_a31_xhdl103;
      wen_a32 <= wen_a32_xhdl104;
      wen_a33 <= wen_a33_xhdl105;
      wen_a34 <= wen_a34_xhdl106;
      wen_a35 <= wen_a35_xhdl107;
      wen_a36 <= wen_a36_xhdl108;
      wen_a37 <= wen_a37_xhdl109;
      wen_a38 <= wen_a38_xhdl110;
      wen_a39 <= wen_a39_xhdl111;
      wen_a40 <= wen_a40_xhdl112;
      wen_a41 <= wen_a41_xhdl113;
      wen_a42 <= wen_a42_xhdl114;
      wen_a43 <= wen_a43_xhdl115;
      wen_a44 <= wen_a44_xhdl116;
      wen_a45 <= wen_a45_xhdl117;
      wen_a46 <= wen_a46_xhdl118;
      wen_a47 <= wen_a47_xhdl119;
      wen_a48 <= wen_a48_xhdl120;
      wen_a49 <= wen_a49_xhdl121;
      wen_a50 <= wen_a50_xhdl122;
      wen_a51 <= wen_a51_xhdl123;
      wen_a52 <= wen_a52_xhdl124;
      wen_a53 <= wen_a53_xhdl125;
      wen_a54 <= wen_a54_xhdl126;
      wen_a55 <= wen_a55_xhdl127;
      wen_a56 <= wen_a56_xhdl128;
      wen_a57 <= wen_a57_xhdl129;
      wen_a58 <= wen_a58_xhdl130;
      wen_a59 <= wen_a59_xhdl131;
      wen_a60 <= wen_a60_xhdl132;
      wen_a61 <= wen_a61_xhdl133;
      wen_a62 <= wen_a62_xhdl134;
      wen_a63 <= wen_a63_xhdl135;
      wen_a64 <= wen_a64_xhdl136;
      wen_a65 <= wen_a65_xhdl137;
      wen_a66 <= wen_a66_xhdl138;
      wen_a67 <= wen_a67_xhdl139;
      wen_a68 <= wen_a68_xhdl140;
      wen_b0 <= wen_b0_xhdl141;
      wen_b1 <= wen_b1_xhdl142;
      wen_b2 <= wen_b2_xhdl143;
      wen_b3 <= wen_b3_xhdl144;
      wen_b4 <= wen_b4_xhdl145;
      wen_b5 <= wen_b5_xhdl146;
      wen_b6 <= wen_b6_xhdl147;
      wen_b7 <= wen_b7_xhdl148;
      wen_b8 <= wen_b8_xhdl149;
      wen_b9 <= wen_b9_xhdl150;
      wen_b10 <= wen_b10_xhdl151;
      wen_b11 <= wen_b11_xhdl152;
      wen_b12 <= wen_b12_xhdl153;
      wen_b13 <= wen_b13_xhdl154;
      wen_b14 <= wen_b14_xhdl155;
      wen_b15 <= wen_b15_xhdl156;
      wen_b16 <= wen_b16_xhdl157;
      wen_b17 <= wen_b17_xhdl158;
      wen_b18 <= wen_b18_xhdl159;
      wen_b19 <= wen_b19_xhdl160;
      wen_b20 <= wen_b20_xhdl161;
      wen_b21 <= wen_b21_xhdl162;
      wen_b22 <= wen_b22_xhdl163;
      wen_b23 <= wen_b23_xhdl164;
      wen_b24 <= wen_b24_xhdl165;
      wen_b25 <= wen_b25_xhdl166;
      wen_b26 <= wen_b26_xhdl167;
      wen_b27 <= wen_b27_xhdl168;
      wen_b28 <= wen_b28_xhdl169;
      wen_b29 <= wen_b29_xhdl170;
      wen_b30 <= wen_b30_xhdl171;
      wen_b31 <= wen_b31_xhdl172;
      wen_b32 <= wen_b32_xhdl173;
      wen_b33 <= wen_b33_xhdl174;
      wen_b34 <= wen_b34_xhdl175;
      wen_b35 <= wen_b35_xhdl176;
      wen_b36 <= wen_b36_xhdl177;
      wen_b37 <= wen_b37_xhdl178;
      wen_b38 <= wen_b38_xhdl179;
      wen_b39 <= wen_b39_xhdl180;
      wen_b40 <= wen_b40_xhdl181;
      wen_b41 <= wen_b41_xhdl182;
      wen_b42 <= wen_b42_xhdl183;
      wen_b43 <= wen_b43_xhdl184;
      wen_b44 <= wen_b44_xhdl185;
      wen_b45 <= wen_b45_xhdl186;
      wen_b46 <= wen_b46_xhdl187;
      wen_b47 <= wen_b47_xhdl188;
      wen_b48 <= wen_b48_xhdl189;
      wen_b49 <= wen_b49_xhdl190;
      wen_b50 <= wen_b50_xhdl191;
      wen_b51 <= wen_b51_xhdl192;
      wen_b52 <= wen_b52_xhdl193;
      wen_b53 <= wen_b53_xhdl194;
      wen_b54 <= wen_b54_xhdl195;
      wen_b55 <= wen_b55_xhdl196;
      wen_b56 <= wen_b56_xhdl197;
      wen_b57 <= wen_b57_xhdl198;
      wen_b58 <= wen_b58_xhdl199;
      wen_b59 <= wen_b59_xhdl200;
      wen_b60 <= wen_b60_xhdl201;
      wen_b61 <= wen_b61_xhdl202;
      wen_b62 <= wen_b62_xhdl203;
      wen_b63 <= wen_b63_xhdl204;
      wen_b64 <= wen_b64_xhdl205;
      wen_b65 <= wen_b65_xhdl206;
      wen_b66 <= wen_b66_xhdl207;
      wen_b67 <= wen_b67_xhdl208;
      wen_b68 <= wen_b68_xhdl209;
      writeData0 <= writeData0_xhdl210;
      writeData1 <= writeData1_xhdl211;
      writeData2 <= writeData2_xhdl212;
      writeData3 <= writeData3_xhdl213;
      writeData4 <= writeData4_xhdl214;
      writeData5 <= writeData5_xhdl215;
      writeData6 <= writeData6_xhdl216;
      writeData7 <= writeData7_xhdl217;
      writeData8 <= writeData8_xhdl218;
      writeData9 <= writeData9_xhdl219;
      writeData10 <= writeData10_xhdl220;
      writeData11 <= writeData11_xhdl221;
      writeData12 <= writeData12_xhdl222;
      writeData13 <= writeData13_xhdl223;
      writeData14 <= writeData14_xhdl224;
      writeData15 <= writeData15_xhdl225;
      writeData16 <= writeData16_xhdl226;
      writeData17 <= writeData17_xhdl227;
      writeData18 <= writeData18_xhdl228;
      writeData19 <= writeData19_xhdl229;
      writeData20 <= writeData20_xhdl230;
      writeData21 <= writeData21_xhdl231;
      writeData22 <= writeData22_xhdl232;
      writeData23 <= writeData23_xhdl233;
      writeData24 <= writeData24_xhdl234;
      writeData25 <= writeData25_xhdl235;
      writeData26 <= writeData26_xhdl236;
      writeData27 <= writeData27_xhdl237;
      writeData28 <= writeData28_xhdl238;
      writeData29 <= writeData29_xhdl239;
      writeData30 <= writeData30_xhdl240;
      writeData31 <= writeData31_xhdl241;
      writeData32 <= writeData32_xhdl242;
      writeData33 <= writeData33_xhdl243;
      writeData34 <= writeData34_xhdl244;
      writeData35 <= writeData35_xhdl245;
      writeData36 <= writeData36_xhdl246;
      writeData37 <= writeData37_xhdl247;
      writeData38 <= writeData38_xhdl248;
      writeData39 <= writeData39_xhdl249;
      writeData40 <= writeData40_xhdl250;
      writeData41 <= writeData41_xhdl251;
      writeData42 <= writeData42_xhdl252;
      writeData43 <= writeData43_xhdl253;
      writeData44 <= writeData44_xhdl254;
      writeData45 <= writeData45_xhdl255;
      writeData46 <= writeData46_xhdl256;
      writeData47 <= writeData47_xhdl257;
      writeData48 <= writeData48_xhdl258;
      writeData49 <= writeData49_xhdl259;
      writeData50 <= writeData50_xhdl260;
      writeData51 <= writeData51_xhdl261;
      writeData52 <= writeData52_xhdl262;
      writeData53 <= writeData53_xhdl263;
      writeData54 <= writeData54_xhdl264;
      writeData55 <= writeData55_xhdl265;
      writeData56 <= writeData56_xhdl266;
      writeData57 <= writeData57_xhdl267;
      writeData58 <= writeData58_xhdl268;
      writeData59 <= writeData59_xhdl269;
      writeData60 <= writeData60_xhdl270;
      writeData61 <= writeData61_xhdl271;
      writeData62 <= writeData62_xhdl272;
      writeData63 <= writeData63_xhdl273;
      writeData64 <= writeData64_xhdl274;
      writeData65 <= writeData65_xhdl275;
      writeData66 <= writeData66_xhdl276;
      writeData67 <= writeData67_xhdl277;
      writeData68 <= writeData68_xhdl278;
      writeAddr0 <= writeAddr0_xhdl279;
      writeAddr1 <= writeAddr1_xhdl280;
      writeAddr2 <= writeAddr2_xhdl281;
      writeAddr3 <= writeAddr3_xhdl282;
      writeAddr4 <= writeAddr4_xhdl283;
      writeAddr5 <= writeAddr5_xhdl284;
      writeAddr6 <= writeAddr6_xhdl285;
      writeAddr7 <= writeAddr7_xhdl286;
      writeAddr8 <= writeAddr8_xhdl287;
      writeAddr9 <= writeAddr9_xhdl288;
      writeAddr10 <= writeAddr10_xhdl289;
      writeAddr11 <= writeAddr11_xhdl290;
      writeAddr12 <= writeAddr12_xhdl291;
      writeAddr13 <= writeAddr13_xhdl292;
      writeAddr14 <= writeAddr14_xhdl293;
      writeAddr15 <= writeAddr15_xhdl294;
      writeAddr16 <= writeAddr16_xhdl295;
      writeAddr17 <= writeAddr17_xhdl296;
      writeAddr18 <= writeAddr18_xhdl297;
      writeAddr19 <= writeAddr19_xhdl298;
      writeAddr20 <= writeAddr20_xhdl299;
      writeAddr21 <= writeAddr21_xhdl300;
      writeAddr22 <= writeAddr22_xhdl301;
      writeAddr23 <= writeAddr23_xhdl302;
      writeAddr24 <= writeAddr24_xhdl303;
      writeAddr25 <= writeAddr25_xhdl304;
      writeAddr26 <= writeAddr26_xhdl305;
      writeAddr27 <= writeAddr27_xhdl306;
      writeAddr28 <= writeAddr28_xhdl307;
      writeAddr29 <= writeAddr29_xhdl308;
      writeAddr30 <= writeAddr30_xhdl309;
      writeAddr31 <= writeAddr31_xhdl310;
      writeAddr32 <= writeAddr32_xhdl311;
      writeAddr33 <= writeAddr33_xhdl312;
      writeAddr34 <= writeAddr34_xhdl313;
      writeAddr35 <= writeAddr35_xhdl314;
      writeAddr36 <= writeAddr36_xhdl315;
      writeAddr37 <= writeAddr37_xhdl316;
      writeAddr38 <= writeAddr38_xhdl317;
      writeAddr39 <= writeAddr39_xhdl318;
      writeAddr40 <= writeAddr40_xhdl319;
      writeAddr41 <= writeAddr41_xhdl320;
      writeAddr42 <= writeAddr42_xhdl321;
      writeAddr43 <= writeAddr43_xhdl322;
      writeAddr44 <= writeAddr44_xhdl323;
      writeAddr45 <= writeAddr45_xhdl324;
      writeAddr46 <= writeAddr46_xhdl325;
      writeAddr47 <= writeAddr47_xhdl326;
      writeAddr48 <= writeAddr48_xhdl327;
      writeAddr49 <= writeAddr49_xhdl328;
      writeAddr50 <= writeAddr50_xhdl329;
      writeAddr51 <= writeAddr51_xhdl330;
      writeAddr52 <= writeAddr52_xhdl331;
      writeAddr53 <= writeAddr53_xhdl332;
      writeAddr54 <= writeAddr54_xhdl333;
      writeAddr55 <= writeAddr55_xhdl334;
      writeAddr56 <= writeAddr56_xhdl335;
      writeAddr57 <= writeAddr57_xhdl336;
      writeAddr58 <= writeAddr58_xhdl337;
      writeAddr59 <= writeAddr59_xhdl338;
      writeAddr60 <= writeAddr60_xhdl339;
      writeAddr61 <= writeAddr61_xhdl340;
      writeAddr62 <= writeAddr62_xhdl341;
      writeAddr63 <= writeAddr63_xhdl342;
      writeAddr64 <= writeAddr64_xhdl343;
      writeAddr65 <= writeAddr65_xhdl344;
      writeAddr66 <= writeAddr66_xhdl345;
      writeAddr67 <= writeAddr67_xhdl346;
      writeAddr68 <= writeAddr68_xhdl347;
      readAddr0 <= readAddr0_xhdl348;
      readAddr1 <= readAddr1_xhdl349;
      readAddr2 <= readAddr2_xhdl350;
      readAddr3 <= readAddr3_xhdl351;
      readAddr4 <= readAddr4_xhdl352;
      readAddr5 <= readAddr5_xhdl353;
      readAddr6 <= readAddr6_xhdl354;
      readAddr7 <= readAddr7_xhdl355;
      readAddr8 <= readAddr8_xhdl356;
      readAddr9 <= readAddr9_xhdl357;
      readAddr10 <= readAddr10_xhdl358;
      readAddr11 <= readAddr11_xhdl359;
      readAddr12 <= readAddr12_xhdl360;
      readAddr13 <= readAddr13_xhdl361;
      readAddr14 <= readAddr14_xhdl362;
      readAddr15 <= readAddr15_xhdl363;
      readAddr16 <= readAddr16_xhdl364;
      readAddr17 <= readAddr17_xhdl365;
      readAddr18 <= readAddr18_xhdl366;
      readAddr19 <= readAddr19_xhdl367;
      readAddr20 <= readAddr20_xhdl368;
      readAddr21 <= readAddr21_xhdl369;
      readAddr22 <= readAddr22_xhdl370;
      readAddr23 <= readAddr23_xhdl371;
      readAddr24 <= readAddr24_xhdl372;
      readAddr25 <= readAddr25_xhdl373;
      readAddr26 <= readAddr26_xhdl374;
      readAddr27 <= readAddr27_xhdl375;
      readAddr28 <= readAddr28_xhdl376;
      readAddr29 <= readAddr29_xhdl377;
      readAddr30 <= readAddr30_xhdl378;
      readAddr31 <= readAddr31_xhdl379;
      readAddr32 <= readAddr32_xhdl380;
      readAddr33 <= readAddr33_xhdl381;
      readAddr34 <= readAddr34_xhdl382;
      readAddr35 <= readAddr35_xhdl383;
      readAddr36 <= readAddr36_xhdl384;
      readAddr37 <= readAddr37_xhdl385;
      readAddr38 <= readAddr38_xhdl386;
      readAddr39 <= readAddr39_xhdl387;
      readAddr40 <= readAddr40_xhdl388;
      readAddr41 <= readAddr41_xhdl389;
      readAddr42 <= readAddr42_xhdl390;
      readAddr43 <= readAddr43_xhdl391;
      readAddr44 <= readAddr44_xhdl392;
      readAddr45 <= readAddr45_xhdl393;
      readAddr46 <= readAddr46_xhdl394;
      readAddr47 <= readAddr47_xhdl395;
      readAddr48 <= readAddr48_xhdl396;
      readAddr49 <= readAddr49_xhdl397;
      readAddr50 <= readAddr50_xhdl398;
      readAddr51 <= readAddr51_xhdl399;
      readAddr52 <= readAddr52_xhdl400;
      readAddr53 <= readAddr53_xhdl401;
      readAddr54 <= readAddr54_xhdl402;
      readAddr55 <= readAddr55_xhdl403;
      readAddr56 <= readAddr56_xhdl404;
      readAddr57 <= readAddr57_xhdl405;
      readAddr58 <= readAddr58_xhdl406;
      readAddr59 <= readAddr59_xhdl407;
      readAddr60 <= readAddr60_xhdl408;
      readAddr61 <= readAddr61_xhdl409;
      readAddr62 <= readAddr62_xhdl410;
      readAddr63 <= readAddr63_xhdl411;
      readAddr64 <= readAddr64_xhdl412;
      readAddr65 <= readAddr65_xhdl413;
      readAddr66 <= readAddr66_xhdl414;
      readAddr67 <= readAddr67_xhdl415;
      readAddr68 <= readAddr68_xhdl416;
      readData_xhdl1 <= readData_xhdl1_xhdl417;
   END PROCESS;
   
   -- always @ (*)
   ------------------------------------------------------------------------------------------
   -- RAM1K18 blocks
   ------------------------------------------------------------------------------------------
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block68 : RAM1K18 
      PORT MAP (
         A_DOUT => readData68,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData68,
         B_DIN => writeData68,
         A_ADDR => writeAddr68,
         B_ADDR => writeAddr68,
         A_WEN => wen_a68,
         B_WEN => wen_b68,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width68,
         B_WIDTH => width68,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_68,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block67 : RAM1K18 
      PORT MAP (
         A_DOUT => readData67,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData67,
         B_DIN => writeData67,
         A_ADDR => writeAddr67,
         B_ADDR => writeAddr67,
         A_WEN => wen_a67,
         B_WEN => wen_b67,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width67,
         B_WIDTH => width67,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_67,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block66 : RAM1K18 
      PORT MAP (
         A_DOUT => readData66,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData66,
         B_DIN => writeData66,
         A_ADDR => writeAddr66,
         B_ADDR => writeAddr66,
         A_WEN => wen_a66,
         B_WEN => wen_b66,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width66,
         B_WIDTH => width66,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_66,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block65 : RAM1K18 
      PORT MAP (
         A_DOUT => readData65,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData65,
         B_DIN => writeData65,
         A_ADDR => writeAddr65,
         B_ADDR => writeAddr65,
         A_WEN => wen_a65,
         B_WEN => wen_b65,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width65,
         B_WIDTH => width65,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_65,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block64 : RAM1K18 
      PORT MAP (
         A_DOUT => readData64,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData64,
         B_DIN => writeData64,
         A_ADDR => writeAddr64,
         B_ADDR => writeAddr64,
         A_WEN => wen_a64,
         B_WEN => wen_b64,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width64,
         B_WIDTH => width64,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_64,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block63 : RAM1K18 
      PORT MAP (
         A_DOUT => readData63,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData63,
         B_DIN => writeData63,
         A_ADDR => writeAddr63,
         B_ADDR => writeAddr63,
         A_WEN => wen_a63,
         B_WEN => wen_b63,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width63,
         B_WIDTH => width63,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_63,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block62 : RAM1K18 
      PORT MAP (
         A_DOUT => readData62,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData62,
         B_DIN => writeData62,
         A_ADDR => writeAddr62,
         B_ADDR => writeAddr62,
         A_WEN => wen_a62,
         B_WEN => wen_b62,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width62,
         B_WIDTH => width62,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_62,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block61 : RAM1K18 
      PORT MAP (
         A_DOUT => readData61,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData61,
         B_DIN => writeData61,
         A_ADDR => writeAddr61,
         B_ADDR => writeAddr61,
         A_WEN => wen_a61,
         B_WEN => wen_b61,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width61,
         B_WIDTH => width61,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_61,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block60 : RAM1K18 
      PORT MAP (
         A_DOUT => readData60,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData60,
         B_DIN => writeData60,
         A_ADDR => writeAddr60,
         B_ADDR => writeAddr60,
         A_WEN => wen_a60,
         B_WEN => wen_b60,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width60,
         B_WIDTH => width60,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_60,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block59 : RAM1K18 
      PORT MAP (
         A_DOUT => readData59,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData59,
         B_DIN => writeData59,
         A_ADDR => writeAddr59,
         B_ADDR => writeAddr59,
         A_WEN => wen_a59,
         B_WEN => wen_b59,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width59,
         B_WIDTH => width59,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_59,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block58 : RAM1K18 
      PORT MAP (
         A_DOUT => readData58,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData58,
         B_DIN => writeData58,
         A_ADDR => writeAddr58,
         B_ADDR => writeAddr58,
         A_WEN => wen_a58,
         B_WEN => wen_b58,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width58,
         B_WIDTH => width58,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_58,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block57 : RAM1K18 
      PORT MAP (
         A_DOUT => readData57,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData57,
         B_DIN => writeData57,
         A_ADDR => writeAddr57,
         B_ADDR => writeAddr57,
         A_WEN => wen_a57,
         B_WEN => wen_b57,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width57,
         B_WIDTH => width57,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_57,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block56 : RAM1K18 
      PORT MAP (
         A_DOUT => readData56,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData56,
         B_DIN => writeData56,
         A_ADDR => writeAddr56,
         B_ADDR => writeAddr56,
         A_WEN => wen_a56,
         B_WEN => wen_b56,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width56,
         B_WIDTH => width56,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_56,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block55 : RAM1K18 
      PORT MAP (
         A_DOUT => readData55,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData55,
         B_DIN => writeData55,
         A_ADDR => writeAddr55,
         B_ADDR => writeAddr55,
         A_WEN => wen_a55,
         B_WEN => wen_b55,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width55,
         B_WIDTH => width55,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_55,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block54 : RAM1K18 
      PORT MAP (
         A_DOUT => readData54,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData54,
         B_DIN => writeData54,
         A_ADDR => writeAddr54,
         B_ADDR => writeAddr54,
         A_WEN => wen_a54,
         B_WEN => wen_b54,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width54,
         B_WIDTH => width54,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_54,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block53 : RAM1K18 
      PORT MAP (
         A_DOUT => readData53,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData53,
         B_DIN => writeData53,
         A_ADDR => writeAddr53,
         B_ADDR => writeAddr53,
         A_WEN => wen_a53,
         B_WEN => wen_b53,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width53,
         B_WIDTH => width53,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_53,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block52 : RAM1K18 
      PORT MAP (
         A_DOUT => readData52,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData52,
         B_DIN => writeData52,
         A_ADDR => writeAddr52,
         B_ADDR => writeAddr52,
         A_WEN => wen_a52,
         B_WEN => wen_b52,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width52,
         B_WIDTH => width52,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_52,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block51 : RAM1K18 
      PORT MAP (
         A_DOUT => readData51,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData51,
         B_DIN => writeData51,
         A_ADDR => writeAddr51,
         B_ADDR => writeAddr51,
         A_WEN => wen_a51,
         B_WEN => wen_b51,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width51,
         B_WIDTH => width51,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_51,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block50 : RAM1K18 
      PORT MAP (
         A_DOUT => readData50,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData50,
         B_DIN => writeData50,
         A_ADDR => writeAddr50,
         B_ADDR => writeAddr50,
         A_WEN => wen_a50,
         B_WEN => wen_b50,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width50,
         B_WIDTH => width50,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_50,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block49 : RAM1K18 
      PORT MAP (
         A_DOUT => readData49,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData49,
         B_DIN => writeData49,
         A_ADDR => writeAddr49,
         B_ADDR => writeAddr49,
         A_WEN => wen_a49,
         B_WEN => wen_b49,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width49,
         B_WIDTH => width49,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_49,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block48 : RAM1K18 
      PORT MAP (
         A_DOUT => readData48,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData48,
         B_DIN => writeData48,
         A_ADDR => writeAddr48,
         B_ADDR => writeAddr48,
         A_WEN => wen_a48,
         B_WEN => wen_b48,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width48,
         B_WIDTH => width48,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_48,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block47 : RAM1K18 
      PORT MAP (
         A_DOUT => readData47,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData47,
         B_DIN => writeData47,
         A_ADDR => writeAddr47,
         B_ADDR => writeAddr47,
         A_WEN => wen_a47,
         B_WEN => wen_b47,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width47,
         B_WIDTH => width47,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_47,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block46 : RAM1K18 
      PORT MAP (
         A_DOUT => readData46,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData46,
         B_DIN => writeData46,
         A_ADDR => writeAddr46,
         B_ADDR => writeAddr46,
         A_WEN => wen_a46,
         B_WEN => wen_b46,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width46,
         B_WIDTH => width46,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_46,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block45 : RAM1K18 
      PORT MAP (
         A_DOUT => readData45,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData45,
         B_DIN => writeData45,
         A_ADDR => writeAddr45,
         B_ADDR => writeAddr45,
         A_WEN => wen_a45,
         B_WEN => wen_b45,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width45,
         B_WIDTH => width45,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_45,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block44 : RAM1K18 
      PORT MAP (
         A_DOUT => readData44,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData44,
         B_DIN => writeData44,
         A_ADDR => writeAddr44,
         B_ADDR => writeAddr44,
         A_WEN => wen_a44,
         B_WEN => wen_b44,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width44,
         B_WIDTH => width44,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_44,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block43 : RAM1K18 
      PORT MAP (
         A_DOUT => readData43,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData43,
         B_DIN => writeData43,
         A_ADDR => writeAddr43,
         B_ADDR => writeAddr43,
         A_WEN => wen_a43,
         B_WEN => wen_b43,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width43,
         B_WIDTH => width43,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_43,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block42 : RAM1K18 
      PORT MAP (
         A_DOUT => readData42,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData42,
         B_DIN => writeData42,
         A_ADDR => writeAddr42,
         B_ADDR => writeAddr42,
         A_WEN => wen_a42,
         B_WEN => wen_b42,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width42,
         B_WIDTH => width42,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_42,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block41 : RAM1K18 
      PORT MAP (
         A_DOUT => readData41,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData41,
         B_DIN => writeData41,
         A_ADDR => writeAddr41,
         B_ADDR => writeAddr41,
         A_WEN => wen_a41,
         B_WEN => wen_b41,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width41,
         B_WIDTH => width41,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_41,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block40 : RAM1K18 
      PORT MAP (
         A_DOUT => readData40,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData40,
         B_DIN => writeData40,
         A_ADDR => writeAddr40,
         B_ADDR => writeAddr40,
         A_WEN => wen_a40,
         B_WEN => wen_b40,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width40,
         B_WIDTH => width40,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_40,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block39 : RAM1K18 
      PORT MAP (
         A_DOUT => readData39,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData39,
         B_DIN => writeData39,
         A_ADDR => writeAddr39,
         B_ADDR => writeAddr39,
         A_WEN => wen_a39,
         B_WEN => wen_b39,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width39,
         B_WIDTH => width39,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_39,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block38 : RAM1K18 
      PORT MAP (
         A_DOUT => readData38,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData38,
         B_DIN => writeData38,
         A_ADDR => writeAddr38,
         B_ADDR => writeAddr38,
         A_WEN => wen_a38,
         B_WEN => wen_b38,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width38,
         B_WIDTH => width38,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_38,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block37 : RAM1K18 
      PORT MAP (
         A_DOUT => readData37,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData37,
         B_DIN => writeData37,
         A_ADDR => writeAddr37,
         B_ADDR => writeAddr37,
         A_WEN => wen_a37,
         B_WEN => wen_b37,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width37,
         B_WIDTH => width37,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_37,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block36 : RAM1K18 
      PORT MAP (
         A_DOUT => readData36,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData36,
         B_DIN => writeData36,
         A_ADDR => writeAddr36,
         B_ADDR => writeAddr36,
         A_WEN => wen_a36,
         B_WEN => wen_b36,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width36,
         B_WIDTH => width36,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_36,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block35 : RAM1K18 
      PORT MAP (
         A_DOUT => readData35,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData35,
         B_DIN => writeData35,
         A_ADDR => writeAddr35,
         B_ADDR => writeAddr35,
         A_WEN => wen_a35,
         B_WEN => wen_b35,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width35,
         B_WIDTH => width35,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_35,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block34 : RAM1K18 
      PORT MAP (
         A_DOUT => readData34,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData34,
         B_DIN => writeData34,
         A_ADDR => writeAddr34,
         B_ADDR => writeAddr34,
         A_WEN => wen_a34,
         B_WEN => wen_b34,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width34,
         B_WIDTH => width34,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_34,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block33 : RAM1K18 
      PORT MAP (
         A_DOUT => readData33,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData33,
         B_DIN => writeData33,
         A_ADDR => writeAddr33,
         B_ADDR => writeAddr33,
         A_WEN => wen_a33,
         B_WEN => wen_b33,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width33,
         B_WIDTH => width33,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_33,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block32 : RAM1K18 
      PORT MAP (
         A_DOUT => readData32,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData32,
         B_DIN => writeData32,
         A_ADDR => writeAddr32,
         B_ADDR => writeAddr32,
         A_WEN => wen_a32,
         B_WEN => wen_b32,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width32,
         B_WIDTH => width32,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_32,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block31 : RAM1K18 
      PORT MAP (
         A_DOUT => readData31,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData31,
         B_DIN => writeData31,
         A_ADDR => writeAddr31,
         B_ADDR => writeAddr31,
         A_WEN => wen_a31,
         B_WEN => wen_b31,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width31,
         B_WIDTH => width31,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_31,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block30 : RAM1K18 
      PORT MAP (
         A_DOUT => readData30,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData30,
         B_DIN => writeData30,
         A_ADDR => writeAddr30,
         B_ADDR => writeAddr30,
         A_WEN => wen_a30,
         B_WEN => wen_b30,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width30,
         B_WIDTH => width30,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_30,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block29 : RAM1K18 
      PORT MAP (
         A_DOUT => readData29,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData29,
         B_DIN => writeData29,
         A_ADDR => writeAddr29,
         B_ADDR => writeAddr29,
         A_WEN => wen_a29,
         B_WEN => wen_b29,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width29,
         B_WIDTH => width29,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_29,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block28 : RAM1K18 
      PORT MAP (
         A_DOUT => readData28,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData28,
         B_DIN => writeData28,
         A_ADDR => writeAddr28,
         B_ADDR => writeAddr28,
         A_WEN => wen_a28,
         B_WEN => wen_b28,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width28,
         B_WIDTH => width28,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_28,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block27 : RAM1K18 
      PORT MAP (
         A_DOUT => readData27,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData27,
         B_DIN => writeData27,
         A_ADDR => writeAddr27,
         B_ADDR => writeAddr27,
         A_WEN => wen_a27,
         B_WEN => wen_b27,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width27,
         B_WIDTH => width27,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_27,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block26 : RAM1K18 
      PORT MAP (
         A_DOUT => readData26,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData26,
         B_DIN => writeData26,
         A_ADDR => writeAddr26,
         B_ADDR => writeAddr26,
         A_WEN => wen_a26,
         B_WEN => wen_b26,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width26,
         B_WIDTH => width26,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_26,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block25 : RAM1K18 
      PORT MAP (
         A_DOUT => readData25,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData25,
         B_DIN => writeData25,
         A_ADDR => writeAddr25,
         B_ADDR => writeAddr25,
         A_WEN => wen_a25,
         B_WEN => wen_b25,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width25,
         B_WIDTH => width25,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_25,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block24 : RAM1K18 
      PORT MAP (
         A_DOUT => readData24,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData24,
         B_DIN => writeData24,
         A_ADDR => writeAddr24,
         B_ADDR => writeAddr24,
         A_WEN => wen_a24,
         B_WEN => wen_b24,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width24,
         B_WIDTH => width24,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_24,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block23 : RAM1K18 
      PORT MAP (
         A_DOUT => readData23,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData23,
         B_DIN => writeData23,
         A_ADDR => writeAddr23,
         B_ADDR => writeAddr23,
         A_WEN => wen_a23,
         B_WEN => wen_b23,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width23,
         B_WIDTH => width23,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_23,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block22 : RAM1K18 
      PORT MAP (
         A_DOUT => readData22,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData22,
         B_DIN => writeData22,
         A_ADDR => writeAddr22,
         B_ADDR => writeAddr22,
         A_WEN => wen_a22,
         B_WEN => wen_b22,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width22,
         B_WIDTH => width22,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_22,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block21 : RAM1K18 
      PORT MAP (
         A_DOUT => readData21,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData21,
         B_DIN => writeData21,
         A_ADDR => writeAddr21,
         B_ADDR => writeAddr21,
         A_WEN => wen_a21,
         B_WEN => wen_b21,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width21,
         B_WIDTH => width21,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_21,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block20 : RAM1K18 
      PORT MAP (
         A_DOUT => readData20,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData20,
         B_DIN => writeData20,
         A_ADDR => writeAddr20,
         B_ADDR => writeAddr20,
         A_WEN => wen_a20,
         B_WEN => wen_b20,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width20,
         B_WIDTH => width20,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_20,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block19 : RAM1K18 
      PORT MAP (
         A_DOUT => readData19,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData19,
         B_DIN => writeData19,
         A_ADDR => writeAddr19,
         B_ADDR => writeAddr19,
         A_WEN => wen_a19,
         B_WEN => wen_b19,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width19,
         B_WIDTH => width19,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_19,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block18 : RAM1K18 
      PORT MAP (
         A_DOUT => readData18,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData18,
         B_DIN => writeData18,
         A_ADDR => writeAddr18,
         B_ADDR => writeAddr18,
         A_WEN => wen_a18,
         B_WEN => wen_b18,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width18,
         B_WIDTH => width18,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_18,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block17 : RAM1K18 
      PORT MAP (
         A_DOUT => readData17,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData17,
         B_DIN => writeData17,
         A_ADDR => writeAddr17,
         B_ADDR => writeAddr17,
         A_WEN => wen_a17,
         B_WEN => wen_b17,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width17,
         B_WIDTH => width17,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_17,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block16 : RAM1K18 
      PORT MAP (
         A_DOUT => readData16,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData16,
         B_DIN => writeData16,
         A_ADDR => writeAddr16,
         B_ADDR => writeAddr16,
         A_WEN => wen_a16,
         B_WEN => wen_b16,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width16,
         B_WIDTH => width16,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_16,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block15 : RAM1K18 
      PORT MAP (
         A_DOUT => readData15,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData15,
         B_DIN => writeData15,
         A_ADDR => writeAddr15,
         B_ADDR => writeAddr15,
         A_WEN => wen_a15,
         B_WEN => wen_b15,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width15,
         B_WIDTH => width15,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_15,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block14 : RAM1K18 
      PORT MAP (
         A_DOUT => readData14,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData14,
         B_DIN => writeData14,
         A_ADDR => writeAddr14,
         B_ADDR => writeAddr14,
         A_WEN => wen_a14,
         B_WEN => wen_b14,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width14,
         B_WIDTH => width14,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_14,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block13 : RAM1K18 
      PORT MAP (
         A_DOUT => readData13,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData13,
         B_DIN => writeData13,
         A_ADDR => writeAddr13,
         B_ADDR => writeAddr13,
         A_WEN => wen_a13,
         B_WEN => wen_b13,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width13,
         B_WIDTH => width13,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_13,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block12 : RAM1K18 
      PORT MAP (
         A_DOUT => readData12,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData12,
         B_DIN => writeData12,
         A_ADDR => writeAddr12,
         B_ADDR => writeAddr12,
         A_WEN => wen_a12,
         B_WEN => wen_b12,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width12,
         B_WIDTH => width12,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_12,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block11 : RAM1K18 
      PORT MAP (
         A_DOUT => readData11,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData11,
         B_DIN => writeData11,
         A_ADDR => writeAddr11,
         B_ADDR => writeAddr11,
         A_WEN => wen_a11,
         B_WEN => wen_b11,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width11,
         B_WIDTH => width11,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_11,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block10 : RAM1K18 
      PORT MAP (
         A_DOUT => readData10,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData10,
         B_DIN => writeData10,
         A_ADDR => writeAddr10,
         B_ADDR => writeAddr10,
         A_WEN => wen_a10,
         B_WEN => wen_b10,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width10,
         B_WIDTH => width10,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_10,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block9 : RAM1K18 
      PORT MAP (
         A_DOUT => readData9,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData9,
         B_DIN => writeData9,
         A_ADDR => writeAddr9,
         B_ADDR => writeAddr9,
         A_WEN => wen_a9,
         B_WEN => wen_b9,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width9,
         B_WIDTH => width9,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_9,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block8 : RAM1K18 
      PORT MAP (
         A_DOUT => readData8,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData8,
         B_DIN => writeData8,
         A_ADDR => writeAddr8,
         B_ADDR => writeAddr8,
         A_WEN => wen_a8,
         B_WEN => wen_b8,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width8,
         B_WIDTH => width8,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_8,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block7 : RAM1K18 
      PORT MAP (
         A_DOUT => readData7,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData7,
         B_DIN => writeData7,
         A_ADDR => writeAddr7,
         B_ADDR => writeAddr7,
         A_WEN => wen_a7,
         B_WEN => wen_b7,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width7,
         B_WIDTH => width7,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_7,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block6 : RAM1K18 
      PORT MAP (
         A_DOUT => readData6,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData6,
         B_DIN => writeData6,
         A_ADDR => writeAddr6,
         B_ADDR => writeAddr6,
         A_WEN => wen_a6,
         B_WEN => wen_b6,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width6,
         B_WIDTH => width6,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_6,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block5 : RAM1K18 
      PORT MAP (
         A_DOUT => readData5,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData5,
         B_DIN => writeData5,
         A_ADDR => writeAddr5,
         B_ADDR => writeAddr5,
         A_WEN => wen_a5,
         B_WEN => wen_b5,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width5,
         B_WIDTH => width5,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_5,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block4 : RAM1K18 
      PORT MAP (
         A_DOUT => readData4,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData4,
         B_DIN => writeData4,
         A_ADDR => writeAddr4,
         B_ADDR => writeAddr4,
         A_WEN => wen_a4,
         B_WEN => wen_b4,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width4,
         B_WIDTH => width4,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_4,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block3 : RAM1K18 
      PORT MAP (
         A_DOUT => readData3,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData3,
         B_DIN => writeData3,
         A_ADDR => writeAddr3,
         B_ADDR => writeAddr3,
         A_WEN => wen_a3,
         B_WEN => wen_b3,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width3,
         B_WIDTH => width3,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_3,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block2 : RAM1K18 
      PORT MAP (
         A_DOUT => readData2,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData2,
         B_DIN => writeData2,
         A_ADDR => writeAddr2,
         B_ADDR => writeAddr2,
         A_WEN => wen_a2,
         B_WEN => wen_b2,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width2,
         B_WIDTH => width2,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_2,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block1 : RAM1K18 
      PORT MAP (
         A_DOUT => readData1,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData1,
         B_DIN => writeData1,
         A_ADDR => writeAddr1,
         B_ADDR => writeAddr1,
         A_WEN => wen_a1,
         B_WEN => wen_b1,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width1,
         B_WIDTH => width1,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_1,
         SII_LOCK => '0');   
   
   -- <<X-HDL>> Can't find translated component 'RAM1K18'. Port & generic names and types may not match. No template will be included
   block0 : RAM1K18 
      PORT MAP (
         A_DOUT => readData0,
         B_DOUT => open,
         A_CLK => clk,
         B_CLK => clk,
         A_ARST_N => resetn,
         B_ARST_N => resetn,
         A_BLK => "111",
         B_BLK => "000",
         A_DIN => writeData0,
         B_DIN => writeData0,
         A_ADDR => writeAddr0,
         B_ADDR => writeAddr0,
         A_WEN => wen_a0,
         B_WEN => wen_b0,
         A_DOUT_CLK => '1',
         B_DOUT_CLK => '1',
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_ARST_N => '1',
         B_DOUT_ARST_N => '1',
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_DOUT_LAT => '1',
         B_DOUT_LAT => '1',
         A_WIDTH => width0,
         B_WIDTH => width0,
         A_WMODE => '0',
         B_WMODE => '0',
         A_EN => '1',
         B_EN => '1',
         BUSY => lsram_2k_BUSY_0,
         SII_LOCK => '0');   
   
   lsram_2k_BUSY_all_xhdl2 <= lsram_2k_BUSY_0 OR lsram_2k_BUSY_1 OR 
   lsram_2k_BUSY_2 OR lsram_2k_BUSY_3 OR lsram_2k_BUSY_4 OR 
   lsram_2k_BUSY_5 OR lsram_2k_BUSY_6 OR lsram_2k_BUSY_7 OR 
   lsram_2k_BUSY_8 OR lsram_2k_BUSY_9 OR lsram_2k_BUSY_10 OR 
   lsram_2k_BUSY_11 OR lsram_2k_BUSY_12 OR lsram_2k_BUSY_13 OR 
   lsram_2k_BUSY_14 OR lsram_2k_BUSY_15 OR lsram_2k_BUSY_16 OR 
   lsram_2k_BUSY_17 OR lsram_2k_BUSY_18 OR lsram_2k_BUSY_19 OR 
   lsram_2k_BUSY_20 OR lsram_2k_BUSY_21 OR lsram_2k_BUSY_22 OR 
   lsram_2k_BUSY_23 OR lsram_2k_BUSY_24 OR lsram_2k_BUSY_25 OR 
   lsram_2k_BUSY_26 OR lsram_2k_BUSY_27 OR lsram_2k_BUSY_28 OR 
   lsram_2k_BUSY_29 OR lsram_2k_BUSY_30 OR lsram_2k_BUSY_31 OR 
   lsram_2k_BUSY_32 OR lsram_2k_BUSY_33 OR lsram_2k_BUSY_34 OR 
   lsram_2k_BUSY_35 OR lsram_2k_BUSY_36 OR lsram_2k_BUSY_37 OR 
   lsram_2k_BUSY_38 OR lsram_2k_BUSY_39 OR lsram_2k_BUSY_40 OR 
   lsram_2k_BUSY_41 OR lsram_2k_BUSY_42 OR lsram_2k_BUSY_43 OR 
   lsram_2k_BUSY_44 OR lsram_2k_BUSY_45 OR lsram_2k_BUSY_46 OR 
   lsram_2k_BUSY_47 OR lsram_2k_BUSY_48 OR lsram_2k_BUSY_49 OR 
   lsram_2k_BUSY_50 OR lsram_2k_BUSY_51 OR lsram_2k_BUSY_52 OR 
   lsram_2k_BUSY_53 OR lsram_2k_BUSY_54 OR lsram_2k_BUSY_55 OR 
   lsram_2k_BUSY_56 OR lsram_2k_BUSY_57 OR lsram_2k_BUSY_58 OR 
   lsram_2k_BUSY_59 OR lsram_2k_BUSY_60 OR lsram_2k_BUSY_61 OR 
   lsram_2k_BUSY_62 OR lsram_2k_BUSY_63 OR lsram_2k_BUSY_64 OR 
   lsram_2k_BUSY_65 OR lsram_2k_BUSY_66 OR lsram_2k_BUSY_67 OR 
   lsram_2k_BUSY_68 ;

END ARCHITECTURE translated;
