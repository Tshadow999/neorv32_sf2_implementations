-- ********************************************************************/
-- Actel Corporation Proprietary and Confidential
--  Copyright 2011 Actel Corporation.  All rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
-- ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
-- IN ADVANCE IN WRITING.
--
-- Description:  SRAM block, 4 byte wide, 64 to 2304 deep (in steps
--               of 64 for Word accesses), 64 to 4608 deep (in steps
--               of 64 for Half-Word accesses) and 64 to 4608 deep (in 
--               steps of 128 for Byte accesses) used to construct 
--               the memory.
--
-- Revision Information:
-- Date     Description
--
-- SVN Revision Information:
-- SVN $Revision: 4805 $
-- SVN $Date: 2008-11-27 17:48:48 +0530 (Thu, 27 Nov 2008) $
--
-- Resolved SARs
-- SAR      Date     Who   Description
--
-- Notes:
--
-- ********************************************************************/
library ieee;
use     ieee.std_logic_1164.all;
use     ieee.std_logic_arith.all;
use     ieee.std_logic_unsigned.all;
use     ieee.std_logic_misc.all;

ENTITY COREAPBLSRAM_C0_COREAPBLSRAM_C0_0_usram_64to4608x16 IS
   GENERIC (
      -- ---------------------------------------------------------------------
      -- Parameters
      -- ---------------------------------------------------------------------
      -- DEPTH can range from
      -- 64 to 4608bytes  , in steps of 64bytes
      USRAM_NUM_LOCATIONS_DWIDTH16   :  integer := 64;    
      APB_DWIDTH                     :  integer := 32);    
   PORT (
      -- ---------------------------------------------------------------------
-- Port declarations
-- ---------------------------------------------------------------------
-- AhbFabric interface
-- Inputs

      writeData               : IN std_logic_vector(APB_DWIDTH - 1 DOWNTO 0);   
      -- Output

      readData                : OUT std_logic_vector(APB_DWIDTH - 1 
      DOWNTO 0);   
-- Inputs

      wen                     : IN std_logic;   
      ren                     : IN std_logic;   
      writeAddr               : IN std_logic_vector(17 DOWNTO 0);   
      readAddr                : IN std_logic_vector(17 DOWNTO 0);   
      clk                     : IN std_logic;   
      resetn                  : IN std_logic;   
      u_4K_BUSY_all              : OUT std_logic);   
END ENTITY COREAPBLSRAM_C0_COREAPBLSRAM_C0_0_usram_64to4608x16;

ARCHITECTURE translated OF COREAPBLSRAM_C0_COREAPBLSRAM_C0_0_usram_64to4608x16 IS

   COMPONENT RAM64x18 
      PORT (
         A_DOUT               : OUT std_logic_vector(17 DOWNTO 0); 
         B_DOUT               : OUT std_logic_vector(17 DOWNTO 0); 
         A_ADDR_CLK                : IN std_logic;
         B_ADDR_CLK                : IN std_logic; 
         A_ADDR_EN              : IN std_logic;
         B_ADDR_EN              : IN std_logic;
         A_ADDR_LAT              : IN std_logic;
         B_ADDR_LAT              : IN std_logic;
         A_ADDR_ARST_N                : IN std_logic; 
         B_ADDR_ARST_N                 : IN std_logic;
         A_ADDR_SRST_N                : IN std_logic; 
         B_ADDR_SRST_N                 : IN std_logic;
         A_DOUT_CLK                : IN std_logic;
         B_DOUT_CLK                : IN std_logic;
         A_DOUT_EN                : IN std_logic;
         B_DOUT_EN                : IN std_logic;
         A_DOUT_LAT                : IN std_logic;
         B_DOUT_LAT                : IN std_logic;
        A_DOUT_ARST_N                : IN std_logic;
         B_DOUT_ARST_N                : IN std_logic;
         A_DOUT_SRST_N                : IN std_logic;
         B_DOUT_SRST_N                : IN std_logic;
         A_ADDR              : IN std_logic_vector(9 DOWNTO 0);
         B_ADDR              : IN std_logic_vector(9 DOWNTO 0);
         A_WIDTH              : IN std_logic_vector(2 DOWNTO 0);
         B_WIDTH              : IN std_logic_vector(2 DOWNTO 0);
         A_BLK              : IN std_logic_vector(1 DOWNTO 0);
         B_BLK              : IN std_logic_vector(1 DOWNTO 0);
         A_EN                : IN std_logic;
         B_EN                : IN std_logic;
         C_CLK                : IN std_logic; 
         C_BLK              : IN std_logic_vector(1 DOWNTO 0);
         C_DIN              : IN std_logic_vector(17 DOWNTO 0);
        C_EN                : IN std_logic;
        C_ADDR              : IN std_logic_vector(9 DOWNTO 0);
         C_WEN              : IN std_logic;
         C_WIDTH              : IN std_logic_vector(2 DOWNTO 0);    
        BUSY                : OUT std_logic;
         SII_LOCK                : IN std_logic);
  END COMPONENT;   

   -- ---------------------------------------------------------------------
   -- Constant declarations
   -- ---------------------------------------------------------------------
   -- ---------------------------------------------------------------------
   -- Signal declarations
   -- ---------------------------------------------------------------------
   SIGNAL ckRdAddr                 :  std_logic_vector(13 DOWNTO 6);   
   SIGNAL width0                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width1                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width2                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width3                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width4                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width5                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width6                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width7                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width8                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width9                   :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width10                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width11                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width12                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width13                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width14                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width15                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width16                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width17                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width18                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width19                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width20                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width21                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width22                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width23                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width24                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width25                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width26                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width27                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width28                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width29                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width30                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width31                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width32                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width33                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width34                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width35                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width36                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width37                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width38                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width39                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width40                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width41                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width42                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width43                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width44                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width45                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width46                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width47                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width48                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width49                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width50                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width51                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width52                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width53                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width54                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width55                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width56                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width57                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width58                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width59                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width60                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width61                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width62                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width63                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width64                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width65                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width66                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width67                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width68                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width69                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width70                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL width71                  :  std_logic_vector(2 DOWNTO 0);   
   SIGNAL wen_a0                   :  std_logic;   
   SIGNAL wen_a1                   :  std_logic;   
   SIGNAL wen_a2                   :  std_logic;   
   SIGNAL wen_a3                   :  std_logic;   
   SIGNAL wen_a4                   :  std_logic;   
   SIGNAL wen_a5                   :  std_logic;   
   SIGNAL wen_a6                   :  std_logic;   
   SIGNAL wen_a7                   :  std_logic;   
   SIGNAL wen_a8                   :  std_logic;   
   SIGNAL wen_a9                   :  std_logic;   
   SIGNAL wen_a10                  :  std_logic;   
   SIGNAL wen_a11                  :  std_logic;   
   SIGNAL wen_a12                  :  std_logic;   
   SIGNAL wen_a13                  :  std_logic;   
   SIGNAL wen_a14                  :  std_logic;   
   SIGNAL wen_a15                  :  std_logic;   
   SIGNAL wen_a16                  :  std_logic;   
   SIGNAL wen_a17                  :  std_logic;   
   SIGNAL wen_a18                  :  std_logic;   
   SIGNAL wen_a19                  :  std_logic;   
   SIGNAL wen_a20                  :  std_logic;   
   SIGNAL wen_a21                  :  std_logic;   
   SIGNAL wen_a22                  :  std_logic;   
   SIGNAL wen_a23                  :  std_logic;   
   SIGNAL wen_a24                  :  std_logic;   
   SIGNAL wen_a25                  :  std_logic;   
   SIGNAL wen_a26                  :  std_logic;   
   SIGNAL wen_a27                  :  std_logic;   
   SIGNAL wen_a28                  :  std_logic;   
   SIGNAL wen_a29                  :  std_logic;   
   SIGNAL wen_a30                  :  std_logic;   
   SIGNAL wen_a31                  :  std_logic;   
   SIGNAL wen_a32                  :  std_logic;   
   SIGNAL wen_a33                  :  std_logic;   
   SIGNAL wen_a34                  :  std_logic;   
   SIGNAL wen_a35                  :  std_logic;   
   SIGNAL wen_a36                  :  std_logic;   
   SIGNAL wen_a37                  :  std_logic;   
   SIGNAL wen_a38                  :  std_logic;   
   SIGNAL wen_a39                  :  std_logic;   
   SIGNAL wen_a40                  :  std_logic;   
   SIGNAL wen_a41                  :  std_logic;   
   SIGNAL wen_a42                  :  std_logic;   
   SIGNAL wen_a43                  :  std_logic;   
   SIGNAL wen_a44                  :  std_logic;   
   SIGNAL wen_a45                  :  std_logic;   
   SIGNAL wen_a46                  :  std_logic;   
   SIGNAL wen_a47                  :  std_logic;   
   SIGNAL wen_a48                  :  std_logic;   
   SIGNAL wen_a49                  :  std_logic;   
   SIGNAL wen_a50                  :  std_logic;   
   SIGNAL wen_a51                  :  std_logic;   
   SIGNAL wen_a52                  :  std_logic;   
   SIGNAL wen_a53                  :  std_logic;   
   SIGNAL wen_a54                  :  std_logic;   
   SIGNAL wen_a55                  :  std_logic;   
   SIGNAL wen_a56                  :  std_logic;   
   SIGNAL wen_a57                  :  std_logic;   
   SIGNAL wen_a58                  :  std_logic;   
   SIGNAL wen_a59                  :  std_logic;   
   SIGNAL wen_a60                  :  std_logic;   
   SIGNAL wen_a61                  :  std_logic;   
   SIGNAL wen_a62                  :  std_logic;   
   SIGNAL wen_a63                  :  std_logic;   
   SIGNAL wen_a64                  :  std_logic;   
   SIGNAL wen_a65                  :  std_logic;   
   SIGNAL wen_a66                  :  std_logic;   
   SIGNAL wen_a67                  :  std_logic;   
   SIGNAL wen_a68                  :  std_logic;   
   SIGNAL wen_a69                  :  std_logic;   
   SIGNAL wen_a70                  :  std_logic;   
   SIGNAL wen_a71                  :  std_logic;   
   SIGNAL wen_b0                   :  std_logic;   
   SIGNAL wen_b1                   :  std_logic;   
   SIGNAL wen_b2                   :  std_logic;   
   SIGNAL wen_b3                   :  std_logic;   
   SIGNAL wen_b4                   :  std_logic;   
   SIGNAL wen_b5                   :  std_logic;   
   SIGNAL wen_b6                   :  std_logic;   
   SIGNAL wen_b7                   :  std_logic;   
   SIGNAL wen_b8                   :  std_logic;   
   SIGNAL wen_b9                   :  std_logic;   
   SIGNAL wen_b10                  :  std_logic;   
   SIGNAL wen_b11                  :  std_logic;   
   SIGNAL wen_b12                  :  std_logic;   
   SIGNAL wen_b13                  :  std_logic;   
   SIGNAL wen_b14                  :  std_logic;   
   SIGNAL wen_b15                  :  std_logic;   
   SIGNAL wen_b16                  :  std_logic;   
   SIGNAL wen_b17                  :  std_logic;   
   SIGNAL wen_b18                  :  std_logic;   
   SIGNAL wen_b19                  :  std_logic;   
   SIGNAL wen_b20                  :  std_logic;   
   SIGNAL wen_b21                  :  std_logic;   
   SIGNAL wen_b22                  :  std_logic;   
   SIGNAL wen_b23                  :  std_logic;   
   SIGNAL wen_b24                  :  std_logic;   
   SIGNAL wen_b25                  :  std_logic;   
   SIGNAL wen_b26                  :  std_logic;   
   SIGNAL wen_b27                  :  std_logic;   
   SIGNAL wen_b28                  :  std_logic;   
   SIGNAL wen_b29                  :  std_logic;   
   SIGNAL wen_b30                  :  std_logic;   
   SIGNAL wen_b31                  :  std_logic;   
   SIGNAL wen_b32                  :  std_logic;   
   SIGNAL wen_b33                  :  std_logic;   
   SIGNAL wen_b34                  :  std_logic;   
   SIGNAL wen_b35                  :  std_logic;   
   SIGNAL wen_b36                  :  std_logic;   
   SIGNAL wen_b37                  :  std_logic;   
   SIGNAL wen_b38                  :  std_logic;   
   SIGNAL wen_b39                  :  std_logic;   
   SIGNAL wen_b40                  :  std_logic;   
   SIGNAL wen_b41                  :  std_logic;   
   SIGNAL wen_b42                  :  std_logic;   
   SIGNAL wen_b43                  :  std_logic;   
   SIGNAL wen_b44                  :  std_logic;   
   SIGNAL wen_b45                  :  std_logic;   
   SIGNAL wen_b46                  :  std_logic;   
   SIGNAL wen_b47                  :  std_logic;   
   SIGNAL wen_b48                  :  std_logic;   
   SIGNAL wen_b49                  :  std_logic;   
   SIGNAL wen_b50                  :  std_logic;   
   SIGNAL wen_b51                  :  std_logic;   
   SIGNAL wen_b52                  :  std_logic;   
   SIGNAL wen_b53                  :  std_logic;   
   SIGNAL wen_b54                  :  std_logic;   
   SIGNAL wen_b55                  :  std_logic;   
   SIGNAL wen_b56                  :  std_logic;   
   SIGNAL wen_b57                  :  std_logic;   
   SIGNAL wen_b58                  :  std_logic;   
   SIGNAL wen_b59                  :  std_logic;   
   SIGNAL wen_b60                  :  std_logic;   
   SIGNAL wen_b61                  :  std_logic;   
   SIGNAL wen_b62                  :  std_logic;   
   SIGNAL wen_b63                  :  std_logic;   
   SIGNAL wen_b64                  :  std_logic;   
   SIGNAL wen_b65                  :  std_logic;   
   SIGNAL wen_b66                  :  std_logic;   
   SIGNAL wen_b67                  :  std_logic;   
   SIGNAL wen_b68                  :  std_logic;   
   SIGNAL wen_b69                  :  std_logic;   
   SIGNAL wen_b70                  :  std_logic;   
   SIGNAL wen_b71                  :  std_logic;   
   SIGNAL writeData0               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData1               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData2               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData3               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData4               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData5               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData6               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData7               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData8               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData9               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData10              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData11              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData12              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData13              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData14              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData15              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData16              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData17              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData18              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData19              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData20              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData21              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData22              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData23              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData24              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData25              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData26              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData27              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData28              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData29              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData30              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData31              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData32              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData33              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData34              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData35              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData36              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData37              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData38              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData39              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData40              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData41              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData42              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData43              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData44              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData45              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData46              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData47              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData48              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData49              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData50              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData51              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData52              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData53              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData54              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData55              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData56              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData57              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData58              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData59              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData60              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData61              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData62              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData63              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData64              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData65              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData66              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData67              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData68              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData69              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData70              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeData71              :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData0                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData1                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData2                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData3                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData4                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData5                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData6                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData7                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData8                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData9                :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData10               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData11               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData12               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData13               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData14               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData15               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData16               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData17               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData18               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData19               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData20               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData21               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData22               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData23               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData24               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData25               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData26               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData27               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData28               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData29               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData30               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData31               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData32               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData33               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData34               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData35               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData36               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData37               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData38               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData39               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData40               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData41               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData42               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData43               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData44               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData45               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData46               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData47               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData48               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData49               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData50               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData51               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData52               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData53               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData54               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData55               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData56               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData57               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData58               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData59               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData60               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData61               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData62               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData63               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData64               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData65               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData66               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData67               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData68               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData69               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData70               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL readData71               :  std_logic_vector(17 DOWNTO 0);   
   SIGNAL writeAddr0               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr1               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr2               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr3               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr4               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr5               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr6               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr7               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr8               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr9               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr10              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr11              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr12              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr13              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr14              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr15              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr16              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr17              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr18              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr19              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr20              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr21              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr22              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr23              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr24              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr25              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr26              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr27              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr28              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr29              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr30              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr31              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr32              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr33              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr34              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr35              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr36              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr37              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr38              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr39              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr40              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr41              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr42              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr43              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr44              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr45              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr46              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr47              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr48              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr49              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr50              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr51              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr52              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr53              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr54              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr55              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr56              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr57              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr58              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr59              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr60              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr61              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr62              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr63              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr64              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr65              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr66              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr67              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr68              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr69              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr70              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL writeAddr71              :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr0                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr1                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr2                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr3                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr4                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr5                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr6                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr7                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr8                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr9                :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr10               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr11               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr12               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr13               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr14               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr15               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr16               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr17               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr18               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr19               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr20               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr21               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr22               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr23               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr24               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr25               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr26               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr27               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr28               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr29               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr30               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr31               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr32               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr33               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr34               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr35               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr36               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr37               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr38               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr39               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr40               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr41               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr42               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr43               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr44               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr45               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr46               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr47               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr48               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr49               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr50               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr51               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr52               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr53               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr54               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr55               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr56               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr57               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr58               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr59               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr60               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr61               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr62               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr63               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr64               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr65               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr66               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr67               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr68               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr69               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr70               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL readAddr71               :  std_logic_vector(9 DOWNTO 0);   
   SIGNAL ablk                     :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL bblk                     :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL cblk                     :  std_logic_vector(1 DOWNTO 0);   
   SIGNAL u_BUSY_71                :  std_logic;   
   SIGNAL u_BUSY_70                :  std_logic;   
   SIGNAL u_BUSY_69                :  std_logic;   
   SIGNAL u_BUSY_68                :  std_logic;   
   SIGNAL u_BUSY_67                :  std_logic;   
   SIGNAL u_BUSY_66                :  std_logic;   
   SIGNAL u_BUSY_65                :  std_logic;   
   SIGNAL u_BUSY_64                :  std_logic;   
   SIGNAL u_BUSY_63                :  std_logic;   
   SIGNAL u_BUSY_62                :  std_logic;   
   SIGNAL u_BUSY_61                :  std_logic;   
   SIGNAL u_BUSY_60                :  std_logic;   
   SIGNAL u_BUSY_59                :  std_logic;   
   SIGNAL u_BUSY_58                :  std_logic;   
   SIGNAL u_BUSY_57                :  std_logic;   
   SIGNAL u_BUSY_56                :  std_logic;   
   SIGNAL u_BUSY_55                :  std_logic;   
   SIGNAL u_BUSY_54                :  std_logic;   
   SIGNAL u_BUSY_53                :  std_logic;   
   SIGNAL u_BUSY_52                :  std_logic;   
   SIGNAL u_BUSY_51                :  std_logic;   
   SIGNAL u_BUSY_50                :  std_logic;   
   SIGNAL u_BUSY_49                :  std_logic;   
   SIGNAL u_BUSY_48                :  std_logic;   
   SIGNAL u_BUSY_47                :  std_logic;   
   SIGNAL u_BUSY_46                :  std_logic;   
   SIGNAL u_BUSY_45                :  std_logic;   
   SIGNAL u_BUSY_44                :  std_logic;   
   SIGNAL u_BUSY_43                :  std_logic;   
   SIGNAL u_BUSY_42                :  std_logic;   
   SIGNAL u_BUSY_41                :  std_logic;   
   SIGNAL u_BUSY_40                :  std_logic;   
   SIGNAL u_BUSY_39                :  std_logic;   
   SIGNAL u_BUSY_38                :  std_logic;   
   SIGNAL u_BUSY_37                :  std_logic;   
   SIGNAL u_BUSY_36                :  std_logic;   
   SIGNAL u_BUSY_35                :  std_logic;   
   SIGNAL u_BUSY_34                :  std_logic;   
   SIGNAL u_BUSY_33                :  std_logic;   
   SIGNAL u_BUSY_32                :  std_logic;   
   SIGNAL u_BUSY_31                :  std_logic;   
   SIGNAL u_BUSY_30                :  std_logic;   
   SIGNAL u_BUSY_29                :  std_logic;   
   SIGNAL u_BUSY_28                :  std_logic;   
   SIGNAL u_BUSY_27                :  std_logic;   
   SIGNAL u_BUSY_26                :  std_logic;   
   SIGNAL u_BUSY_25                :  std_logic;   
   SIGNAL u_BUSY_24                :  std_logic;   
   SIGNAL u_BUSY_23                :  std_logic;   
   SIGNAL u_BUSY_22                :  std_logic;   
   SIGNAL u_BUSY_21                :  std_logic;   
   SIGNAL u_BUSY_20                :  std_logic;   
   SIGNAL u_BUSY_19                :  std_logic;   
   SIGNAL u_BUSY_18                :  std_logic;   
   SIGNAL u_BUSY_17                :  std_logic;   
   SIGNAL u_BUSY_16                :  std_logic;   
   SIGNAL u_BUSY_15                :  std_logic;   
   SIGNAL u_BUSY_14                :  std_logic;   
   SIGNAL u_BUSY_13                :  std_logic;   
   SIGNAL u_BUSY_12                :  std_logic;   
   SIGNAL u_BUSY_11                :  std_logic;   
   SIGNAL u_BUSY_10                :  std_logic;   
   SIGNAL u_BUSY_9                 :  std_logic;   
   SIGNAL u_BUSY_8                 :  std_logic;   
   SIGNAL u_BUSY_7                 :  std_logic;   
   SIGNAL u_BUSY_6                 :  std_logic;   
   SIGNAL u_BUSY_5                 :  std_logic;   
   SIGNAL u_BUSY_4                 :  std_logic;   
   SIGNAL u_BUSY_3                 :  std_logic;   
   SIGNAL u_BUSY_2                 :  std_logic;   
   SIGNAL u_BUSY_1                 :  std_logic;   
   SIGNAL u_BUSY_0                 :  std_logic;   
   SIGNAL readData_xhdl1           :  std_logic_vector(APB_DWIDTH - 1 
   DOWNTO 0);   
   SIGNAL u_4K_BUSY_all_xhdl2         :  std_logic;   

BEGIN
   readData <= readData_xhdl1;
   u_4K_BUSY_all <= u_4K_BUSY_all_xhdl2;

   ------------------------------------------------------------------------
   -- Main body of code
   ------------------------------------------------------------------------
   
   PROCESS (clk, resetn)
   BEGIN
      IF (NOT resetn = '1') THEN
         ckRdAddr(13 DOWNTO 6) <= "00000000";    
      ELSIF (clk'EVENT AND clk = '1') THEN
         ckRdAddr(13 DOWNTO 6) <= readAddr(13 DOWNTO 6);    
      END IF;
   END PROCESS;

   ------------------------------------------------------------------------------------------
   -- Assign values to various signals based on DEPTH and RAM64x16_WIDTH settings.
   -- Default is to build the (byte wide) memory from RAM blocks which are configured to
   -- be tall and narrow.
   ------------------------------------------------------------------------------------------
   
   PROCESS (readData20, readData21, readData22, readData23, readData24, 
   readData25, readData26, readData27, readData60, readData61, 
   readData28, readData62, readData29, 
   readData63, readData64, readData65, readData66, readData67, 
   readData68, readData69, readData30, readData31, writeData, 
   readData32, readData33, readData34, readData35, readData36, 
   readData70, readData37, readData71, 
   readData38, readData39, wen_a0, wen_a1, wen_a2, wen_a3, wen_a4, 
   wen_a5, ckRdAddr, readData40, readData41, readData42, 
   readData43, readData44, readData45, 
   readAddr, readData46, readData47, readData48, readData49, readData10, 
   readData11, readData12, readData13, readData14, readData15, wen, 
   readData16, readData17, readData0, readData50, readData18, readData1, 
   readData51, readData2, readData52, readData19, readData3, 
   readData53, readData4, readData54, 
   readData5, readData6, readData55, readData7, readData56, readData8, 
   readData57, readData9, readData58, readData59, writeAddr)
      VARIABLE width0_xhdl3  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width1_xhdl4  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width2_xhdl5  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width3_xhdl6  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width4_xhdl7  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width5_xhdl8  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width6_xhdl9  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width7_xhdl10  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width8_xhdl11  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width9_xhdl12  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width10_xhdl13  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width11_xhdl14  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width12_xhdl15  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width13_xhdl16  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width14_xhdl17  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width15_xhdl18  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width16_xhdl19  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width17_xhdl20  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width18_xhdl21  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width19_xhdl22  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width20_xhdl23  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width21_xhdl24  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width22_xhdl25  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width23_xhdl26  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width24_xhdl27  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width25_xhdl28  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width26_xhdl29  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width27_xhdl30  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width28_xhdl31  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width29_xhdl32  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width30_xhdl33  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width31_xhdl34  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width32_xhdl35  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width33_xhdl36  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width34_xhdl37  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width35_xhdl38  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width36_xhdl39  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width37_xhdl40  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width38_xhdl41  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width39_xhdl42  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width40_xhdl43  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width41_xhdl44  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width42_xhdl45  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width43_xhdl46  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width44_xhdl47  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width45_xhdl48  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width46_xhdl49  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width47_xhdl50  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width48_xhdl51  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width49_xhdl52  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width50_xhdl53  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width51_xhdl54  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width52_xhdl55  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width53_xhdl56  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width54_xhdl57  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width55_xhdl58  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width56_xhdl59  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width57_xhdl60  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width58_xhdl61  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width59_xhdl62  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width60_xhdl63  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width61_xhdl64  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width62_xhdl65  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width63_xhdl66  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width64_xhdl67  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width65_xhdl68  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width66_xhdl69  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width67_xhdl70  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width68_xhdl71  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width69_xhdl72  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width70_xhdl73  : std_logic_vector(2 DOWNTO 0);
      VARIABLE width71_xhdl74  : std_logic_vector(2 DOWNTO 0);
      VARIABLE wen_a0_xhdl75  : std_logic;
      VARIABLE wen_a1_xhdl76  : std_logic;
      VARIABLE wen_a2_xhdl77  : std_logic;
      VARIABLE wen_a3_xhdl78  : std_logic;
      VARIABLE wen_a4_xhdl79  : std_logic;
      VARIABLE wen_a5_xhdl80  : std_logic;
      VARIABLE wen_a6_xhdl81  : std_logic;
      VARIABLE wen_a7_xhdl82  : std_logic;
      VARIABLE wen_a8_xhdl83  : std_logic;
      VARIABLE wen_a9_xhdl84  : std_logic;
      VARIABLE wen_a10_xhdl85  : std_logic;
      VARIABLE wen_a11_xhdl86  : std_logic;
      VARIABLE wen_a12_xhdl87  : std_logic;
      VARIABLE wen_a13_xhdl88  : std_logic;
      VARIABLE wen_a14_xhdl89  : std_logic;
      VARIABLE wen_a15_xhdl90  : std_logic;
      VARIABLE wen_a16_xhdl91  : std_logic;
      VARIABLE wen_a17_xhdl92  : std_logic;
      VARIABLE wen_a18_xhdl93  : std_logic;
      VARIABLE wen_a19_xhdl94  : std_logic;
      VARIABLE wen_a20_xhdl95  : std_logic;
      VARIABLE wen_a21_xhdl96  : std_logic;
      VARIABLE wen_a22_xhdl97  : std_logic;
      VARIABLE wen_a23_xhdl98  : std_logic;
      VARIABLE wen_a24_xhdl99  : std_logic;
      VARIABLE wen_a25_xhdl100  : std_logic;
      VARIABLE wen_a26_xhdl101  : std_logic;
      VARIABLE wen_a27_xhdl102  : std_logic;
      VARIABLE wen_a28_xhdl103  : std_logic;
      VARIABLE wen_a29_xhdl104  : std_logic;
      VARIABLE wen_a30_xhdl105  : std_logic;
      VARIABLE wen_a31_xhdl106  : std_logic;
      VARIABLE wen_a32_xhdl107  : std_logic;
      VARIABLE wen_a33_xhdl108  : std_logic;
      VARIABLE wen_a34_xhdl109  : std_logic;
      VARIABLE wen_a35_xhdl110  : std_logic;
      VARIABLE wen_a36_xhdl111  : std_logic;
      VARIABLE wen_a37_xhdl112  : std_logic;
      VARIABLE wen_a38_xhdl113  : std_logic;
      VARIABLE wen_a39_xhdl114  : std_logic;
      VARIABLE wen_a40_xhdl115  : std_logic;
      VARIABLE wen_a41_xhdl116  : std_logic;
      VARIABLE wen_a42_xhdl117  : std_logic;
      VARIABLE wen_a43_xhdl118  : std_logic;
      VARIABLE wen_a44_xhdl119  : std_logic;
      VARIABLE wen_a45_xhdl120  : std_logic;
      VARIABLE wen_a46_xhdl121  : std_logic;
      VARIABLE wen_a47_xhdl122  : std_logic;
      VARIABLE wen_a48_xhdl123  : std_logic;
      VARIABLE wen_a49_xhdl124  : std_logic;
      VARIABLE wen_a50_xhdl125  : std_logic;
      VARIABLE wen_a51_xhdl126  : std_logic;
      VARIABLE wen_a52_xhdl127  : std_logic;
      VARIABLE wen_a53_xhdl128  : std_logic;
      VARIABLE wen_a54_xhdl129  : std_logic;
      VARIABLE wen_a55_xhdl130  : std_logic;
      VARIABLE wen_a56_xhdl131  : std_logic;
      VARIABLE wen_a57_xhdl132  : std_logic;
      VARIABLE wen_a58_xhdl133  : std_logic;
      VARIABLE wen_a59_xhdl134  : std_logic;
      VARIABLE wen_a60_xhdl135  : std_logic;
      VARIABLE wen_a61_xhdl136  : std_logic;
      VARIABLE wen_a62_xhdl137  : std_logic;
      VARIABLE wen_a63_xhdl138  : std_logic;
      VARIABLE wen_a64_xhdl139  : std_logic;
      VARIABLE wen_a65_xhdl140  : std_logic;
      VARIABLE wen_a66_xhdl141  : std_logic;
      VARIABLE wen_a67_xhdl142  : std_logic;
      VARIABLE wen_a68_xhdl143  : std_logic;
      VARIABLE wen_a69_xhdl144  : std_logic;
      VARIABLE wen_a70_xhdl145  : std_logic;
      VARIABLE wen_a71_xhdl146  : std_logic;
      VARIABLE wen_b0_xhdl147  : std_logic;
      VARIABLE wen_b1_xhdl148  : std_logic;
      VARIABLE wen_b2_xhdl149  : std_logic;
      VARIABLE wen_b3_xhdl150  : std_logic;
      VARIABLE wen_b4_xhdl151  : std_logic;
      VARIABLE wen_b5_xhdl152  : std_logic;
      VARIABLE wen_b6_xhdl153  : std_logic;
      VARIABLE wen_b7_xhdl154  : std_logic;
      VARIABLE wen_b8_xhdl155  : std_logic;
      VARIABLE wen_b9_xhdl156  : std_logic;
      VARIABLE wen_b10_xhdl157  : std_logic;
      VARIABLE wen_b11_xhdl158  : std_logic;
      VARIABLE wen_b12_xhdl159  : std_logic;
      VARIABLE wen_b13_xhdl160  : std_logic;
      VARIABLE wen_b14_xhdl161  : std_logic;
      VARIABLE wen_b15_xhdl162  : std_logic;
      VARIABLE wen_b16_xhdl163  : std_logic;
      VARIABLE wen_b17_xhdl164  : std_logic;
      VARIABLE wen_b18_xhdl165  : std_logic;
      VARIABLE wen_b19_xhdl166  : std_logic;
      VARIABLE wen_b20_xhdl167  : std_logic;
      VARIABLE wen_b21_xhdl168  : std_logic;
      VARIABLE wen_b22_xhdl169  : std_logic;
      VARIABLE wen_b23_xhdl170  : std_logic;
      VARIABLE wen_b24_xhdl171  : std_logic;
      VARIABLE wen_b25_xhdl172  : std_logic;
      VARIABLE wen_b26_xhdl173  : std_logic;
      VARIABLE wen_b27_xhdl174  : std_logic;
      VARIABLE wen_b28_xhdl175  : std_logic;
      VARIABLE wen_b29_xhdl176  : std_logic;
      VARIABLE wen_b30_xhdl177  : std_logic;
      VARIABLE wen_b31_xhdl178  : std_logic;
      VARIABLE wen_b32_xhdl179  : std_logic;
      VARIABLE wen_b33_xhdl180  : std_logic;
      VARIABLE wen_b34_xhdl181  : std_logic;
      VARIABLE wen_b35_xhdl182  : std_logic;
      VARIABLE wen_b36_xhdl183  : std_logic;
      VARIABLE wen_b37_xhdl184  : std_logic;
      VARIABLE wen_b38_xhdl185  : std_logic;
      VARIABLE wen_b39_xhdl186  : std_logic;
      VARIABLE wen_b40_xhdl187  : std_logic;
      VARIABLE wen_b41_xhdl188  : std_logic;
      VARIABLE wen_b42_xhdl189  : std_logic;
      VARIABLE wen_b43_xhdl190  : std_logic;
      VARIABLE wen_b44_xhdl191  : std_logic;
      VARIABLE wen_b45_xhdl192  : std_logic;
      VARIABLE wen_b46_xhdl193  : std_logic;
      VARIABLE wen_b47_xhdl194  : std_logic;
      VARIABLE wen_b48_xhdl195  : std_logic;
      VARIABLE wen_b49_xhdl196  : std_logic;
      VARIABLE wen_b50_xhdl197  : std_logic;
      VARIABLE wen_b51_xhdl198  : std_logic;
      VARIABLE wen_b52_xhdl199  : std_logic;
      VARIABLE wen_b53_xhdl200  : std_logic;
      VARIABLE wen_b54_xhdl201  : std_logic;
      VARIABLE wen_b55_xhdl202  : std_logic;
      VARIABLE wen_b56_xhdl203  : std_logic;
      VARIABLE wen_b57_xhdl204  : std_logic;
      VARIABLE wen_b58_xhdl205  : std_logic;
      VARIABLE wen_b59_xhdl206  : std_logic;
      VARIABLE wen_b60_xhdl207  : std_logic;
      VARIABLE wen_b61_xhdl208  : std_logic;
      VARIABLE wen_b62_xhdl209  : std_logic;
      VARIABLE wen_b63_xhdl210  : std_logic;
      VARIABLE wen_b64_xhdl211  : std_logic;
      VARIABLE wen_b65_xhdl212  : std_logic;
      VARIABLE wen_b66_xhdl213  : std_logic;
      VARIABLE wen_b67_xhdl214  : std_logic;
      VARIABLE wen_b68_xhdl215  : std_logic;
      VARIABLE wen_b69_xhdl216  : std_logic;
      VARIABLE wen_b70_xhdl217  : std_logic;
      VARIABLE wen_b71_xhdl218  : std_logic;
      VARIABLE writeData0_xhdl219  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData1_xhdl220  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData2_xhdl221  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData3_xhdl222  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData4_xhdl223  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData5_xhdl224  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData6_xhdl225  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData7_xhdl226  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData8_xhdl227  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData9_xhdl228  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData10_xhdl229  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData11_xhdl230  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData12_xhdl231  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData13_xhdl232  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData14_xhdl233  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData15_xhdl234  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData16_xhdl235  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData17_xhdl236  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData18_xhdl237  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData19_xhdl238  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData20_xhdl239  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData21_xhdl240  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData22_xhdl241  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData23_xhdl242  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData24_xhdl243  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData25_xhdl244  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData26_xhdl245  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData27_xhdl246  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData28_xhdl247  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData29_xhdl248  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData30_xhdl249  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData31_xhdl250  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData32_xhdl251  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData33_xhdl252  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData34_xhdl253  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData35_xhdl254  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData36_xhdl255  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData37_xhdl256  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData38_xhdl257  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData39_xhdl258  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData40_xhdl259  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData41_xhdl260  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData42_xhdl261  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData43_xhdl262  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData44_xhdl263  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData45_xhdl264  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData46_xhdl265  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData47_xhdl266  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData48_xhdl267  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData49_xhdl268  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData50_xhdl269  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData51_xhdl270  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData52_xhdl271  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData53_xhdl272  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData54_xhdl273  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData55_xhdl274  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData56_xhdl275  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData57_xhdl276  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData58_xhdl277  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData59_xhdl278  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData60_xhdl279  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData61_xhdl280  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData62_xhdl281  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData63_xhdl282  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData64_xhdl283  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData65_xhdl284  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData66_xhdl285  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData67_xhdl286  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData68_xhdl287  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData69_xhdl288  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData70_xhdl289  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeData71_xhdl290  : std_logic_vector(17 DOWNTO 0);
      VARIABLE writeAddr0_xhdl291  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr1_xhdl292  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr2_xhdl293  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr3_xhdl294  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr4_xhdl295  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr5_xhdl296  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr6_xhdl297  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr7_xhdl298  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr8_xhdl299  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr9_xhdl300  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr10_xhdl301  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr11_xhdl302  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr12_xhdl303  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr13_xhdl304  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr14_xhdl305  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr15_xhdl306  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr16_xhdl307  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr17_xhdl308  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr18_xhdl309  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr19_xhdl310  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr20_xhdl311  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr21_xhdl312  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr22_xhdl313  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr23_xhdl314  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr24_xhdl315  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr25_xhdl316  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr26_xhdl317  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr27_xhdl318  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr28_xhdl319  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr29_xhdl320  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr30_xhdl321  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr31_xhdl322  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr32_xhdl323  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr33_xhdl324  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr34_xhdl325  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr35_xhdl326  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr36_xhdl327  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr37_xhdl328  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr38_xhdl329  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr39_xhdl330  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr40_xhdl331  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr41_xhdl332  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr42_xhdl333  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr43_xhdl334  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr44_xhdl335  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr45_xhdl336  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr46_xhdl337  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr47_xhdl338  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr48_xhdl339  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr49_xhdl340  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr50_xhdl341  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr51_xhdl342  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr52_xhdl343  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr53_xhdl344  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr54_xhdl345  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr55_xhdl346  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr56_xhdl347  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr57_xhdl348  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr58_xhdl349  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr59_xhdl350  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr60_xhdl351  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr61_xhdl352  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr62_xhdl353  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr63_xhdl354  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr64_xhdl355  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr65_xhdl356  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr66_xhdl357  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr67_xhdl358  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr68_xhdl359  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr69_xhdl360  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr70_xhdl361  : std_logic_vector(9 DOWNTO 0);
      VARIABLE writeAddr71_xhdl362  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr0_xhdl363  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr1_xhdl364  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr2_xhdl365  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr3_xhdl366  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr4_xhdl367  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr5_xhdl368  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr6_xhdl369  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr7_xhdl370  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr8_xhdl371  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr9_xhdl372  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr10_xhdl373  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr11_xhdl374  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr12_xhdl375  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr13_xhdl376  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr14_xhdl377  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr15_xhdl378  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr16_xhdl379  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr17_xhdl380  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr18_xhdl381  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr19_xhdl382  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr20_xhdl383  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr21_xhdl384  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr22_xhdl385  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr23_xhdl386  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr24_xhdl387  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr25_xhdl388  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr26_xhdl389  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr27_xhdl390  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr28_xhdl391  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr29_xhdl392  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr30_xhdl393  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr31_xhdl394  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr32_xhdl395  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr33_xhdl396  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr34_xhdl397  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr35_xhdl398  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr36_xhdl399  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr37_xhdl400  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr38_xhdl401  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr39_xhdl402  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr40_xhdl403  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr41_xhdl404  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr42_xhdl405  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr43_xhdl406  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr44_xhdl407  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr45_xhdl408  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr46_xhdl409  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr47_xhdl410  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr48_xhdl411  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr49_xhdl412  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr50_xhdl413  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr51_xhdl414  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr52_xhdl415  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr53_xhdl416  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr54_xhdl417  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr55_xhdl418  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr56_xhdl419  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr57_xhdl420  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr58_xhdl421  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr59_xhdl422  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr60_xhdl423  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr61_xhdl424  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr62_xhdl425  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr63_xhdl426  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr64_xhdl427  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr65_xhdl428  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr66_xhdl429  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr67_xhdl430  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr68_xhdl431  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr69_xhdl432  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr70_xhdl433  : std_logic_vector(9 DOWNTO 0);
      VARIABLE readAddr71_xhdl434  : std_logic_vector(9 DOWNTO 0);
      VARIABLE ablk_xhdl435  : std_logic_vector(1 DOWNTO 0);
      VARIABLE bblk_xhdl436  : std_logic_vector(1 DOWNTO 0);
      VARIABLE cblk_xhdl437  : std_logic_vector(1 DOWNTO 0);
      VARIABLE readData_xhdl1_xhdl437_w16  : std_logic_vector(15
      DOWNTO 0);
      
      VARIABLE xhdl438  : std_logic_vector(5 DOWNTO 0);
      VARIABLE xhdl439  : std_logic_vector(2 DOWNTO 0);
   BEGIN
      width0_xhdl3 := "000";    
      width1_xhdl4 := "000";    
      width2_xhdl5 := "000";    
      width3_xhdl6 := "000";    
      width4_xhdl7 := "000";    
      width5_xhdl8 := "000";    
      width6_xhdl9 := "000";    
      width7_xhdl10 := "000";    
      width8_xhdl11 := "000";    
      width9_xhdl12 := "000";    
      width10_xhdl13 := "000";    
      width11_xhdl14 := "000";    
      width12_xhdl15 := "000";    
      width13_xhdl16 := "000";    
      width14_xhdl17 := "000";    
      width15_xhdl18 := "000";    
      width16_xhdl19 := "000";    
      width17_xhdl20 := "000";    
      width18_xhdl21 := "000";    
      width19_xhdl22 := "000";    
      width20_xhdl23 := "000";    
      width21_xhdl24 := "000";    
      width22_xhdl25 := "000";    
      width23_xhdl26 := "000";    
      width24_xhdl27 := "000";    
      width25_xhdl28 := "000";    
      width26_xhdl29 := "000";    
      width27_xhdl30 := "000";    
      width28_xhdl31 := "000";    
      width29_xhdl32 := "000";    
      width30_xhdl33 := "000";    
      width31_xhdl34 := "000";    
      width32_xhdl35 := "000";    
      width33_xhdl36 := "000";    
      width34_xhdl37 := "000";    
      width35_xhdl38 := "000";    
      width36_xhdl39 := "000";    
      width37_xhdl40 := "000";    
      width38_xhdl41 := "000";    
      width39_xhdl42 := "000";    
      width40_xhdl43 := "000";    
      width41_xhdl44 := "000";    
      width42_xhdl45 := "000";    
      width43_xhdl46 := "000";    
      width44_xhdl47 := "000";    
      width45_xhdl48 := "000";    
      width46_xhdl49 := "000";    
      width47_xhdl50 := "000";    
      width48_xhdl51 := "000";    
      width49_xhdl52 := "000";    
      width50_xhdl53 := "000";    
      width51_xhdl54 := "000";    
      width52_xhdl55 := "000";    
      width53_xhdl56 := "000";    
      width54_xhdl57 := "000";    
      width55_xhdl58 := "000";    
      width56_xhdl59 := "000";    
      width57_xhdl60 := "000";    
      width58_xhdl61 := "000";    
      width59_xhdl62 := "000";    
      width60_xhdl63 := "000";    
      width61_xhdl64 := "000";    
      width62_xhdl65 := "000";    
      width63_xhdl66 := "000";    
      width64_xhdl67 := "000";    
      width65_xhdl68 := "000";    
      width66_xhdl69 := "000";    
      width67_xhdl70 := "000";    
      width68_xhdl71 := "000";    
      width69_xhdl72 := "000";    
      width70_xhdl73 := "000";    
      width71_xhdl74 := "000";    
      wen_a0_xhdl75 := '0';    
      wen_a1_xhdl76 := '0';    
      wen_a2_xhdl77 := '0';    
      wen_a3_xhdl78 := '0';    
      wen_a4_xhdl79 := '0';    
      wen_a5_xhdl80 := '0';    
      wen_a6_xhdl81 := '0';    
      wen_a7_xhdl82 := '0';    
      wen_a8_xhdl83 := '0';    
      wen_a9_xhdl84 := '0';    
      wen_a10_xhdl85 := '0';    
      wen_a11_xhdl86 := '0';    
      wen_a12_xhdl87 := '0';    
      wen_a13_xhdl88 := '0';    
      wen_a14_xhdl89 := '0';    
      wen_a15_xhdl90 := '0';    
      wen_a16_xhdl91 := '0';    
      wen_a17_xhdl92 := '0';    
      wen_a18_xhdl93 := '0';    
      wen_a19_xhdl94 := '0';    
      wen_a20_xhdl95 := '0';    
      wen_a21_xhdl96 := '0';    
      wen_a22_xhdl97 := '0';    
      wen_a23_xhdl98 := '0';    
      wen_a24_xhdl99 := '0';    
      wen_a25_xhdl100 := '0';    
      wen_a26_xhdl101 := '0';    
      wen_a27_xhdl102 := '0';    
      wen_a28_xhdl103 := '0';    
      wen_a29_xhdl104 := '0';    
      wen_a30_xhdl105 := '0';    
      wen_a31_xhdl106 := '0';    
      wen_a32_xhdl107 := '0';    
      wen_a33_xhdl108 := '0';    
      wen_a34_xhdl109 := '0';    
      wen_a35_xhdl110 := '0';    
      wen_a36_xhdl111 := '0';    
      wen_a37_xhdl112 := '0';    
      wen_a38_xhdl113 := '0';    
      wen_a39_xhdl114 := '0';    
      wen_a40_xhdl115 := '0';    
      wen_a41_xhdl116 := '0';    
      wen_a42_xhdl117 := '0';    
      wen_a43_xhdl118 := '0';    
      wen_a44_xhdl119 := '0';    
      wen_a45_xhdl120 := '0';    
      wen_a46_xhdl121 := '0';    
      wen_a47_xhdl122 := '0';    
      wen_a48_xhdl123 := '0';    
      wen_a49_xhdl124 := '0';    
      wen_a50_xhdl125 := '0';    
      wen_a51_xhdl126 := '0';    
      wen_a52_xhdl127 := '0';    
      wen_a53_xhdl128 := '0';    
      wen_a54_xhdl129 := '0';    
      wen_a55_xhdl130 := '0';    
      wen_a56_xhdl131 := '0';    
      wen_a57_xhdl132 := '0';    
      wen_a58_xhdl133 := '0';    
      wen_a59_xhdl134 := '0';    
      wen_a60_xhdl135 := '0';    
      wen_a61_xhdl136 := '0';    
      wen_a62_xhdl137 := '0';    
      wen_a63_xhdl138 := '0';    
      wen_a64_xhdl139 := '0';    
      wen_a65_xhdl140 := '0';    
      wen_a66_xhdl141 := '0';    
      wen_a67_xhdl142 := '0';    
      wen_a68_xhdl143 := '0';    
      wen_a69_xhdl144 := '0';    
      wen_a70_xhdl145 := '0';    
      wen_a71_xhdl146 := '0';    
      wen_b0_xhdl147 := '0';    
      wen_b1_xhdl148 := '0';    
      wen_b2_xhdl149 := '0';    
      wen_b3_xhdl150 := '0';    
      wen_b4_xhdl151 := '0';    
      wen_b5_xhdl152 := '0';    
      wen_b6_xhdl153 := '0';    
      wen_b7_xhdl154 := '0';    
      wen_b8_xhdl155 := '0';    
      wen_b9_xhdl156 := '0';    
      wen_b10_xhdl157 := '0';    
      wen_b11_xhdl158 := '0';    
      wen_b12_xhdl159 := '0';    
      wen_b13_xhdl160 := '0';    
      wen_b14_xhdl161 := '0';    
      wen_b15_xhdl162 := '0';    
      wen_b16_xhdl163 := '0';    
      wen_b17_xhdl164 := '0';    
      wen_b18_xhdl165 := '0';    
      wen_b19_xhdl166 := '0';    
      wen_b20_xhdl167 := '0';    
      wen_b21_xhdl168 := '0';    
      wen_b22_xhdl169 := '0';    
      wen_b23_xhdl170 := '0';    
      wen_b24_xhdl171 := '0';    
      wen_b25_xhdl172 := '0';    
      wen_b26_xhdl173 := '0';    
      wen_b27_xhdl174 := '0';    
      wen_b28_xhdl175 := '0';    
      wen_b29_xhdl176 := '0';    
      wen_b30_xhdl177 := '0';    
      wen_b31_xhdl178 := '0';    
      wen_b32_xhdl179 := '0';    
      wen_b33_xhdl180 := '0';    
      wen_b34_xhdl181 := '0';    
      wen_b35_xhdl182 := '0';    
      wen_b36_xhdl183 := '0';    
      wen_b37_xhdl184 := '0';    
      wen_b38_xhdl185 := '0';    
      wen_b39_xhdl186 := '0';    
      wen_b40_xhdl187 := '0';    
      wen_b41_xhdl188 := '0';    
      wen_b42_xhdl189 := '0';    
      wen_b43_xhdl190 := '0';    
      wen_b44_xhdl191 := '0';    
      wen_b45_xhdl192 := '0';    
      wen_b46_xhdl193 := '0';    
      wen_b47_xhdl194 := '0';    
      wen_b48_xhdl195 := '0';    
      wen_b49_xhdl196 := '0';    
      wen_b50_xhdl197 := '0';    
      wen_b51_xhdl198 := '0';    
      wen_b52_xhdl199 := '0';    
      wen_b53_xhdl200 := '0';    
      wen_b54_xhdl201 := '0';    
      wen_b55_xhdl202 := '0';    
      wen_b56_xhdl203 := '0';    
      wen_b57_xhdl204 := '0';    
      wen_b58_xhdl205 := '0';    
      wen_b59_xhdl206 := '0';    
      wen_b60_xhdl207 := '0';    
      wen_b61_xhdl208 := '0';    
      wen_b62_xhdl209 := '0';    
      wen_b63_xhdl210 := '0';    
      wen_b64_xhdl211 := '0';    
      wen_b65_xhdl212 := '0';    
      wen_b66_xhdl213 := '0';    
      wen_b67_xhdl214 := '0';    
      wen_b68_xhdl215 := '0';    
      wen_b69_xhdl216 := '0';    
      wen_b70_xhdl217 := '0';    
      wen_b71_xhdl218 := '0';    
      writeData0_xhdl219 := "000000000000000000";    
      writeData1_xhdl220 := "000000000000000000";    
      writeData2_xhdl221 := "000000000000000000";    
      writeData3_xhdl222 := "000000000000000000";    
      writeData4_xhdl223 := "000000000000000000";    
      writeData5_xhdl224 := "000000000000000000";    
      writeData6_xhdl225 := "000000000000000000";    
      writeData7_xhdl226 := "000000000000000000";    
      writeData8_xhdl227 := "000000000000000000";    
      writeData9_xhdl228 := "000000000000000000";    
      writeData10_xhdl229 := "000000000000000000";    
      writeData11_xhdl230 := "000000000000000000";    
      writeData12_xhdl231 := "000000000000000000";    
      writeData13_xhdl232 := "000000000000000000";    
      writeData14_xhdl233 := "000000000000000000";    
      writeData15_xhdl234 := "000000000000000000";    
      writeData16_xhdl235 := "000000000000000000";    
      writeData17_xhdl236 := "000000000000000000";    
      writeData18_xhdl237 := "000000000000000000";    
      writeData19_xhdl238 := "000000000000000000";    
      writeData20_xhdl239 := "000000000000000000";    
      writeData21_xhdl240 := "000000000000000000";    
      writeData22_xhdl241 := "000000000000000000";    
      writeData23_xhdl242 := "000000000000000000";    
      writeData24_xhdl243 := "000000000000000000";    
      writeData25_xhdl244 := "000000000000000000";    
      writeData26_xhdl245 := "000000000000000000";    
      writeData27_xhdl246 := "000000000000000000";    
      writeData28_xhdl247 := "000000000000000000";    
      writeData29_xhdl248 := "000000000000000000";    
      writeData30_xhdl249 := "000000000000000000";    
      writeData31_xhdl250 := "000000000000000000";    
      writeData32_xhdl251 := "000000000000000000";    
      writeData33_xhdl252 := "000000000000000000";    
      writeData34_xhdl253 := "000000000000000000";    
      writeData35_xhdl254 := "000000000000000000";    
      writeData36_xhdl255 := "000000000000000000";    
      writeData37_xhdl256 := "000000000000000000";    
      writeData38_xhdl257 := "000000000000000000";    
      writeData39_xhdl258 := "000000000000000000";    
      writeData40_xhdl259 := "000000000000000000";    
      writeData41_xhdl260 := "000000000000000000";    
      writeData42_xhdl261 := "000000000000000000";    
      writeData43_xhdl262 := "000000000000000000";    
      writeData44_xhdl263 := "000000000000000000";    
      writeData45_xhdl264 := "000000000000000000";    
      writeData46_xhdl265 := "000000000000000000";    
      writeData47_xhdl266 := "000000000000000000";    
      writeData48_xhdl267 := "000000000000000000";    
      writeData49_xhdl268 := "000000000000000000";    
      writeData50_xhdl269 := "000000000000000000";    
      writeData51_xhdl270 := "000000000000000000";    
      writeData52_xhdl271 := "000000000000000000";    
      writeData53_xhdl272 := "000000000000000000";    
      writeData54_xhdl273 := "000000000000000000";    
      writeData55_xhdl274 := "000000000000000000";    
      writeData56_xhdl275 := "000000000000000000";    
      writeData57_xhdl276 := "000000000000000000";    
      writeData58_xhdl277 := "000000000000000000";    
      writeData59_xhdl278 := "000000000000000000";    
      writeData60_xhdl279 := "000000000000000000";    
      writeData61_xhdl280 := "000000000000000000";    
      writeData62_xhdl281 := "000000000000000000";    
      writeData63_xhdl282 := "000000000000000000";    
      writeData64_xhdl283 := "000000000000000000";    
      writeData65_xhdl284 := "000000000000000000";    
      writeData66_xhdl285 := "000000000000000000";    
      writeData67_xhdl286 := "000000000000000000";    
      writeData68_xhdl287 := "000000000000000000";    
      writeData69_xhdl288 := "000000000000000000";    
      writeData70_xhdl289 := "000000000000000000";    
      writeData71_xhdl290 := "000000000000000000";    
      writeAddr0_xhdl291 := "0000000000";    
      writeAddr1_xhdl292 := "0000000000";    
      writeAddr2_xhdl293 := "0000000000";    
      writeAddr3_xhdl294 := "0000000000";    
      writeAddr4_xhdl295 := "0000000000";    
      writeAddr5_xhdl296 := "0000000000";    
      writeAddr6_xhdl297 := "0000000000";    
      writeAddr7_xhdl298 := "0000000000";    
      writeAddr8_xhdl299 := "0000000000";    
      writeAddr9_xhdl300 := "0000000000";    
      writeAddr10_xhdl301 := "0000000000";    
      writeAddr11_xhdl302 := "0000000000";    
      writeAddr12_xhdl303 := "0000000000";    
      writeAddr13_xhdl304 := "0000000000";    
      writeAddr14_xhdl305 := "0000000000";    
      writeAddr15_xhdl306 := "0000000000";    
      writeAddr16_xhdl307 := "0000000000";    
      writeAddr17_xhdl308 := "0000000000";    
      writeAddr18_xhdl309 := "0000000000";    
      writeAddr19_xhdl310 := "0000000000";    
      writeAddr20_xhdl311 := "0000000000";    
      writeAddr21_xhdl312 := "0000000000";    
      writeAddr22_xhdl313 := "0000000000";    
      writeAddr23_xhdl314 := "0000000000";    
      writeAddr24_xhdl315 := "0000000000";    
      writeAddr25_xhdl316 := "0000000000";    
      writeAddr26_xhdl317 := "0000000000";    
      writeAddr27_xhdl318 := "0000000000";    
      writeAddr28_xhdl319 := "0000000000";    
      writeAddr29_xhdl320 := "0000000000";    
      writeAddr30_xhdl321 := "0000000000";    
      writeAddr31_xhdl322 := "0000000000";    
      writeAddr32_xhdl323 := "0000000000";    
      writeAddr33_xhdl324 := "0000000000";    
      writeAddr34_xhdl325 := "0000000000";    
      writeAddr35_xhdl326 := "0000000000";    
      writeAddr36_xhdl327 := "0000000000";    
      writeAddr37_xhdl328 := "0000000000";    
      writeAddr38_xhdl329 := "0000000000";    
      writeAddr39_xhdl330 := "0000000000";    
      writeAddr40_xhdl331 := "0000000000";    
      writeAddr41_xhdl332 := "0000000000";    
      writeAddr42_xhdl333 := "0000000000";    
      writeAddr43_xhdl334 := "0000000000";    
      writeAddr44_xhdl335 := "0000000000";    
      writeAddr45_xhdl336 := "0000000000";    
      writeAddr46_xhdl337 := "0000000000";    
      writeAddr47_xhdl338 := "0000000000";    
      writeAddr48_xhdl339 := "0000000000";    
      writeAddr49_xhdl340 := "0000000000";    
      writeAddr50_xhdl341 := "0000000000";    
      writeAddr51_xhdl342 := "0000000000";    
      writeAddr52_xhdl343 := "0000000000";    
      writeAddr53_xhdl344 := "0000000000";    
      writeAddr54_xhdl345 := "0000000000";    
      writeAddr55_xhdl346 := "0000000000";    
      writeAddr56_xhdl347 := "0000000000";    
      writeAddr57_xhdl348 := "0000000000";    
      writeAddr58_xhdl349 := "0000000000";    
      writeAddr59_xhdl350 := "0000000000";    
      writeAddr60_xhdl351 := "0000000000";    
      writeAddr61_xhdl352 := "0000000000";    
      writeAddr62_xhdl353 := "0000000000";    
      writeAddr63_xhdl354 := "0000000000";    
      writeAddr64_xhdl355 := "0000000000";    
      writeAddr65_xhdl356 := "0000000000";    
      writeAddr66_xhdl357 := "0000000000";    
      writeAddr67_xhdl358 := "0000000000";    
      writeAddr68_xhdl359 := "0000000000";    
      writeAddr69_xhdl360 := "0000000000";    
      writeAddr70_xhdl361 := "0000000000";    
      writeAddr71_xhdl362 := "0000000000";    
      readAddr0_xhdl363 := "0000000000";    
      readAddr1_xhdl364 := "0000000000";    
      readAddr2_xhdl365 := "0000000000";    
      readAddr3_xhdl366 := "0000000000";    
      readAddr4_xhdl367 := "0000000000";    
      readAddr5_xhdl368 := "0000000000";    
      readAddr6_xhdl369 := "0000000000";    
      readAddr7_xhdl370 := "0000000000";    
      readAddr8_xhdl371 := "0000000000";    
      readAddr9_xhdl372 := "0000000000";    
      readAddr10_xhdl373 := "0000000000";    
      readAddr11_xhdl374 := "0000000000";    
      readAddr12_xhdl375 := "0000000000";    
      readAddr13_xhdl376 := "0000000000";    
      readAddr14_xhdl377 := "0000000000";    
      readAddr15_xhdl378 := "0000000000";    
      readAddr16_xhdl379 := "0000000000";    
      readAddr17_xhdl380 := "0000000000";    
      readAddr18_xhdl381 := "0000000000";    
      readAddr19_xhdl382 := "0000000000";    
      readAddr20_xhdl383 := "0000000000";    
      readAddr21_xhdl384 := "0000000000";    
      readAddr22_xhdl385 := "0000000000";    
      readAddr23_xhdl386 := "0000000000";    
      readAddr24_xhdl387 := "0000000000";    
      readAddr25_xhdl388 := "0000000000";    
      readAddr26_xhdl389 := "0000000000";    
      readAddr27_xhdl390 := "0000000000";    
      readAddr28_xhdl391 := "0000000000";    
      readAddr29_xhdl392 := "0000000000";    
      readAddr30_xhdl393 := "0000000000";    
      readAddr31_xhdl394 := "0000000000";    
      readAddr32_xhdl395 := "0000000000";    
      readAddr33_xhdl396 := "0000000000";    
      readAddr34_xhdl397 := "0000000000";    
      readAddr35_xhdl398 := "0000000000";    
      readAddr36_xhdl399 := "0000000000";    
      readAddr37_xhdl400 := "0000000000";    
      readAddr38_xhdl401 := "0000000000";    
      readAddr39_xhdl402 := "0000000000";    
      readAddr40_xhdl403 := "0000000000";    
      readAddr41_xhdl404 := "0000000000";    
      readAddr42_xhdl405 := "0000000000";    
      readAddr43_xhdl406 := "0000000000";    
      readAddr44_xhdl407 := "0000000000";    
      readAddr45_xhdl408 := "0000000000";    
      readAddr46_xhdl409 := "0000000000";    
      readAddr47_xhdl410 := "0000000000";    
      readAddr48_xhdl411 := "0000000000";    
      readAddr49_xhdl412 := "0000000000";    
      readAddr50_xhdl413 := "0000000000";    
      readAddr51_xhdl414 := "0000000000";    
      readAddr52_xhdl415 := "0000000000";    
      readAddr53_xhdl416 := "0000000000";    
      readAddr54_xhdl417 := "0000000000";    
      readAddr55_xhdl418 := "0000000000";    
      readAddr56_xhdl419 := "0000000000";    
      readAddr57_xhdl420 := "0000000000";    
      readAddr58_xhdl421 := "0000000000";    
      readAddr59_xhdl422 := "0000000000";    
      readAddr60_xhdl423 := "0000000000";    
      readAddr61_xhdl424 := "0000000000";    
      readAddr62_xhdl425 := "0000000000";    
      readAddr63_xhdl426 := "0000000000";    
      readAddr64_xhdl427 := "0000000000";    
      readAddr65_xhdl428 := "0000000000";    
      readAddr66_xhdl429 := "0000000000";    
      readAddr67_xhdl430 := "0000000000";    
      readAddr68_xhdl431 := "0000000000";    
      readAddr69_xhdl432 := "0000000000";    
      readAddr70_xhdl433 := "0000000000";    
      readAddr71_xhdl434 := "0000000000";    
      ablk_xhdl435 := "00";    
      bblk_xhdl436 := "00";
        
            IF (APB_DWIDTH = 16) THEN
               
               --ablk_xhdl435 := "11";    
               --bblk_xhdl436 := "11";    
               ablk_xhdl435 := ren & ren;    
               bblk_xhdl436 := ren & ren;
               cblk_xhdl437 := wen & wen;
               CASE USRAM_NUM_LOCATIONS_DWIDTH16 IS
                  WHEN 64 =>
                           -- RAM 0 and RAM 1 for 64x32 configuration
                           
                           width0_xhdl3 := "100";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           wen_a0_xhdl75 := wen;    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           readData_xhdl1_xhdl437_w16 := readData0(16 DOWNTO 9) & readData0(7 DOWNTO 
                           0);    
                  WHEN 128 =>
                           -- RAM 1 to RAM 4 for 64x32 configuration
                           
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           wen_a2_xhdl77 := wen;    
                           wen_a1_xhdl76 := wen;    
                           readData_xhdl1_xhdl437_w16 := readData2(7 DOWNTO 0) & readData1(7 DOWNTO 
                           0);    
                  WHEN 192 =>
                           -- RAM 0 to RAM 5 for 64x32 configuration
                           
                           width3_xhdl6 := "011";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "100";    
                           writeAddr3_xhdl294 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr3_xhdl366 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData3_xhdl222 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData1_xhdl220 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(7 DOWNTO 6) IS
                              WHEN "00" |
                                   "01" =>
                                       --xhdl439 := wen & wen & '0';  
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';  				       
                              WHEN "10" =>
                                       --xhdl439 := '0' & '0' & wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;  				       
                              WHEN OTHERS  =>
                                       --xhdl439 := '0' & '0' & '0';  
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';  				       
                              
                           END CASE;
                           CASE ckRdAddr(7 DOWNTO 6) IS
                              WHEN "00" |
                                   "01" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData3(7 DOWNTO 0) & readData2(7 DOWNTO 0)
                                       ;    
                              WHEN "10" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData1(16 
                                       DOWNTO 9) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 256 =>
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           wen_a4_xhdl79 := wen;    
                           wen_a3_xhdl78 := wen;    
                           wen_a2_xhdl77 := wen;    
                           wen_a1_xhdl76 := wen;    
                           readData_xhdl1_xhdl437_w16 := 
                           readData4(3 DOWNTO 0) & readData3(3 DOWNTO 
                           0) & readData2(3 DOWNTO 0) & readData1(3 
                           DOWNTO 0);    
                  WHEN 320 =>
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "100";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(8 DOWNTO 6) IS
                              WHEN "000" |
                                   "001" |
                                   "010" |
                                   "011" =>
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                              WHEN "100" =>
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                              WHEN OTHERS  =>
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(8 DOWNTO 6) IS
                              WHEN "000" |
                                   "001" |
                                   "010" |
                                   "011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData1(16 
                                       DOWNTO 9) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 384 =>
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(8 DOWNTO 6) IS
                              WHEN "000" |
                                   "001" |
                                   "010" |
                                   "011" =>
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100" |
                                   "101" =>
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(8 DOWNTO 6) IS
                              WHEN "000" |
                                   "001" |
                                   "010" |
                                   "011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "100" |
                                   "101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 448 =>
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(8 DOWNTO 6) IS
                              WHEN "000" |
                                   "001" |
                                   "010" |
                                   "011" =>
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100" |
                                   "101" =>
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110" =>
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(8 DOWNTO 6) IS
                              WHEN "000" |
                                   "001" |
                                   "010" |
                                   "011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "100" |
                                   "101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData2(7 DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 512 =>
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           wen_a8_xhdl83 := wen;    
                           wen_a7_xhdl82 := wen;    
                           wen_a6_xhdl81 := wen;    
                           wen_a5_xhdl80 := wen;    
                           wen_a4_xhdl79 := wen;    
                           wen_a3_xhdl78 := wen;    
                           wen_a2_xhdl77 := wen;    
                           wen_a1_xhdl76 := wen;    
                           readData_xhdl1_xhdl437_w16 := readData8(1 DOWNTO 0) & readData7(1 DOWNTO 0) & 
			   readData6(1 DOWNTO 0) & readData5(1 DOWNTO 0) & readData4(1 DOWNTO 0) & 
                           readData3(1 DOWNTO 0) & readData2(1 DOWNTO 0) 
                           & readData1(1 DOWNTO 0);    
                  WHEN 576 =>
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "100";    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" =>
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData8(1 DOWNTO 0) & readData7(1 DOWNTO 0) 
                                       & readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0);    
                              WHEN "1000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData0(16 DOWNTO 9) & readData0(7 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 640 =>
                           --512x2   
                           
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           -- 128x8
                           
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" |
                                   "1001" =>
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                       readData9(1 DOWNTO 0) & readData8(1 DOWNTO 0) 
                                       & readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0);    
                              WHEN "1000" |
                                   "1001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 704 =>
                           --512x2   
                           
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" |
                                   "1001" =>
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1010" =>
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData10(1 
                                       DOWNTO 0) & readData9(1 DOWNTO 0) 
                                       & readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0);    
                              WHEN "1000" |
                                   "1001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "1010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 768 =>
                           --512x2   
                           
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData11(1 
                                       DOWNTO 0) & readData10(1 DOWNTO 0)
                                       & readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0);    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 832 =>
                           --512x2
                           
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1100" =>
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData12(1 
                                       DOWNTO 0) & readData11(1 DOWNTO 0)
                                       & readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0);    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "1100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 896 =>
                           --512x2
                           
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1100" |
                                   "1101" =>
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData13(1 
                                       DOWNTO 0) & readData12(1 DOWNTO 0)
                                       & readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0);    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "1100" |
                                   "1101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 960 =>
                           --512x2
                           
                           width14_xhdl17 := "001";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr14_xhdl305 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr14_xhdl377 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData14_xhdl233 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1100" |
                                   "1101" =>
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1110" =>
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(9 DOWNTO 6) IS
                              WHEN "0000" |
                                   "0001" |
                                   "0010" |
                                   "0011" |
                                   "0100" |
                                   "0101" |
                                   "0110" |
                                   "0111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData14(1 
                                       DOWNTO 0) & readData13(1 DOWNTO 0)
                                       & readData12(1 DOWNTO 0) & 
                                       readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0);    
                              WHEN "1000" |
                                   "1001" |
                                   "1010" |
                                   "1011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "1100" |
                                   "1101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "1110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1024 =>
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "000";    
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(9 DOWNTO 0);  
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(9 DOWNTO 0);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(15);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(14);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(13);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(12);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(11);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(10);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(9);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(8);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(7);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(6);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(5);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(4);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(3);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(2);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(1);    
                           writeData0_xhdl219 := "00000000000000000" & 
                           writeData(0);    
                           wen_a15_xhdl90 := wen;    
                           wen_a14_xhdl89 := wen;    
                           wen_a13_xhdl88 := wen;    
                           wen_a12_xhdl87 := wen;    
                           wen_a11_xhdl86 := wen;    
                           wen_a10_xhdl85 := wen;    
                           wen_a9_xhdl84 := wen;    
                           wen_a8_xhdl83 := wen;    
                           wen_a7_xhdl82 := wen;    
                           wen_a6_xhdl81 := wen;    
                           wen_a5_xhdl80 := wen;    
                           wen_a4_xhdl79 := wen;    
                           wen_a3_xhdl78 := wen;    
                           wen_a2_xhdl77 := wen;    
                           wen_a1_xhdl76 := wen;    
                           wen_a0_xhdl75 := wen;    
                           readData_xhdl1_xhdl437_w16 := readData15(0) & readData14(0) & 
                           readData13(0) & readData12(0) & readData11(0) 
                           & readData10(0) & readData9(0) & readData8(0) 
                           & readData7(0) & readData6(0) & readData5(0) 
                           & readData4(0) & readData3(0) & readData2(0) 
                           & readData1(0) & readData0(0);    
                  WHEN 1088 =>
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "100";    
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(15);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(14);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(13);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(12);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(11);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(10);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(9);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(8);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(7);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(6);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(5);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(4);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(3);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(2);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(1);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" =>
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData16(0)
                                       & readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0) & readData2(0) & 
                                       readData1(0);    
                              WHEN "10000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1152 =>
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(15);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(14);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(13);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(12);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(11);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(10);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(9);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(8);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(7);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(6);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(5);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(4);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(3);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(2);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(1);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" =>
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData17(0)
                                       & readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0);    
                              WHEN "10000" |
                                   "10001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1216 =>
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(15);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(14);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(13);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(12);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(11);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(10);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(9);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(8);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(7);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(6);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(5);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(4);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(3);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(2);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(1);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" =>
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10010" =>
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData18(0)
                                       & readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0);    
                              WHEN "10000" |
                                   "10001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "10010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1280 =>
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(15);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(14);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(13);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(12);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(11);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(10);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(9);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(8);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(7);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(6);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(5);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(4);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(3);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(2);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(1);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData19(0)
                                       & readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1344 =>
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(15);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(14);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(13);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(12);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(11);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(10);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(9);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(8);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(7);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(6);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(5);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(4);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(3);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(2);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(1);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10100" =>
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData20(0)
                                       & readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "10100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1408 =>
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(15);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(14);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(13);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(12);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(11);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(10);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(9);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(8);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(7);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(6);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(5);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(4);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(3);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(2);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(1);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10100" |
                                   "10101" =>
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData21(0)
                                       & readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "10100" |
                                   "10101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1472 =>
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(15);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(14);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(13);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(12);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(11);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(10);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(9);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(8);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(7);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(6);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(5);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(4);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(3);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(2);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(1);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10100" |
                                   "10101" =>
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10110" =>
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData22(0)
                                       & readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "10100" |
                                   "10101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "10110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1536 =>
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "001";    
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(15);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(14);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(13);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(12);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(11);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(10);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(9);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(8);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(7);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(6);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(5);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(4);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(3);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(2);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(1);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(0);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData0_xhdl219 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData23(0)
                                       & readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData7(1 
                                       DOWNTO 0) & readData6(1 DOWNTO 0) 
                                       & readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0) & 
                                       readData0(1 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1600 =>
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "100";    
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(15);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(14);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(13);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(12);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(11);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(10);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(9);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(8);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(7);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(6);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(5);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(4);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(3);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(2);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(1);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(0);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" =>
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData24(0)
                                       & readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData8(1 
                                       DOWNTO 0) & readData7(1 DOWNTO 0) 
                                       & readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0);    
                              WHEN "11000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1664 =>
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(15);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(14);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(13);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(12);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(11);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(10);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(9);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(8);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(7);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(6);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(5);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(4);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(3);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(2);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(1);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(0);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" |
                                   "11001" =>
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData25(0)
                                       & readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData9(1 
                                       DOWNTO 0) & readData8(1 DOWNTO 0) 
                                       & readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0);    
                              WHEN "11000" |
                                   "11001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1728 =>
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(15);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(14);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(13);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(12);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(11);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(10);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(9);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(8);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(7);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(6);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(5);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(4);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(3);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(2);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(1);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(0);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" |
                                   "11001" =>
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11010" =>
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData26(0)
                                       & readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData10(1 
                                       DOWNTO 0) & readData9(1 DOWNTO 0) 
                                       & readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0);    
                              WHEN "11000" |
                                   "11001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "11010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1792 =>
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(15);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(14);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(13);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(12);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(11);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(10);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(9);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(8);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(7);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(6);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(5);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(4);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(3);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(2);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(1);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(0);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData27(0)
                                       & readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData11(1 
                                       DOWNTO 0) & readData10(1 DOWNTO 0)
                                       & readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0);    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1856 =>
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(15);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(14);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(13);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(12);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(11);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(10);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(9);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(8);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(7);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(6);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(5);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(4);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(3);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(2);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(1);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(0);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11100" =>
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData28(0)
                                       & readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData12(1 
                                       DOWNTO 0) & readData11(1 DOWNTO 0)
                                       & readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0);    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "11100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1920 =>
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(15);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(14);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(13);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(12);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(11);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(10);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(9);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(8);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(7);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(6);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(5);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(4);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(3);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(2);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(1);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(0);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11100" |
                                   "11101" =>
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData29(0)
                                       & readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData13(1 
                                       DOWNTO 0) & readData12(1 DOWNTO 0)
                                       & readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0);    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "11100" |
                                   "11101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 1984 =>
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "001";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(15);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(14);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(13);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(12);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(11);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(10);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(9);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(8);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(7);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(6);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(5);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(4);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(3);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(2);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(1);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(0);    
                           writeData14_xhdl233 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11100" |
                                   "11101" =>
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "11110" =>
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                           END CASE;
                           CASE ckRdAddr(10 DOWNTO 6) IS
                              WHEN "00000" |
                                   "00001" |
                                   "00010" |
                                   "00011" |
                                   "00100" |
                                   "00101" |
                                   "00110" |
                                   "00111" |
                                   "01000" |
                                   "01001" |
                                   "01010" |
                                   "01011" |
                                   "01100" |
                                   "01101" |
                                   "01110" |
                                   "01111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData30(0)
                                       & readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0);    
                              WHEN "10000" |
                                   "10001" |
                                   "10010" |
                                   "10011" |
                                   "10100" |
                                   "10101" |
                                   "10110" |
                                   "10111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData14(1 
                                       DOWNTO 0) & readData13(1 DOWNTO 0)
                                       & readData12(1 DOWNTO 0) & 
                                       readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0);    
                              WHEN "11000" |
                                   "11001" |
                                   "11010" |
                                   "11011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "11100" |
                                   "11101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "11110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2048 =>
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "000";    
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(9 DOWNTO 0);  
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(9 DOWNTO 0);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(15);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(14);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(13);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(12);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(11);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(10);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(9);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(8);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(7);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(6);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(5);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(4);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(3);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(2);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(1);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(0);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(15);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(14);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(13);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(12);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(11);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(10);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(9);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(8);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(7);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(6);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(5);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(4);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(3);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(2);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(1);    
                           writeData0_xhdl219 := "00000000000000000" & 
                           writeData(0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData31(0)
                                       & readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData15(0)
                                       & readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0) & readData1(0) & 
                                       readData0(0);    
                              WHEN -- case: 6'b010000, 6'b010001, 6'b010010, 6'b010011, 6'b010100, 6'b010101,6'b010110, 6'b010111, 6'b011000, 6'b011001,...
                              
                              OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                           -- case (ckRdAddr[10:6])
                           
                           
                  WHEN 2112 =>
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "100";    
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(15);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(14);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(13);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(12);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(11);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(10);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(9);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(8);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(7);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(6);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(5);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(4);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(3);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(2);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(1);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(0);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(15);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(14);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(13);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(12);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(11);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(10);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(9);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(8);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(7);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(6);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(5);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(4);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(3);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(2);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(1);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" =>
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData32(0)
                                       & readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData16(0)
                                       & readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0) & readData2(0) & 
                                       readData1(0);    
                              WHEN "100000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2176 =>
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(15);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(14);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(13);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(12);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(11);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(10);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(9);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(8);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(7);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(6);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(5);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(4);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(3);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(2);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(1);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(0);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(15);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(14);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(13);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(12);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(11);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(10);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(9);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(8);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(7);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(6);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(5);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(4);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(3);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(2);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(1);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" =>
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData33(0)
                                       & readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData17(0)
                                       & readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0);    
                              WHEN "100000" |
                                   "100001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2240 =>
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(15);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(14);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(13);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(12);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(11);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(10);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(9);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(8);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(7);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(6);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(5);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(4);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(3);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(2);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(1);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(0);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(15);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(14);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(13);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(12);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(11);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(10);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(9);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(8);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(7);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(6);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(5);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(4);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(3);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(2);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(1);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" =>
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100010" =>
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData34(0)
                                       & readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData18(0)
                                       & readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0);    
                              WHEN "100000" |
                                   "100001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "100010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2304 =>
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(15);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(14);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(13);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(12);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(11);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(10);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(9);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(8);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(7);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(6);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(5);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(4);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(3);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(2);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(1);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(0);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(15);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(14);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(13);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(12);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(11);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(10);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(9);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(8);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(7);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(6);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(5);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(4);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(3);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(2);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(1);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData35(0)
                                       & readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData19(0)
                                       & readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2368 =>
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(15);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(14);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(13);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(12);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(11);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(10);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(9);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(8);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(7);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(6);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(5);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(4);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(3);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(2);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(1);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(0);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(15);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(14);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(13);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(12);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(11);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(10);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(9);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(8);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(7);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(6);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(5);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(4);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(3);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(2);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(1);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100100" =>
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData36(0)
                                       & readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData20(0)
                                       & readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "100100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2432 =>
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(15);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(14);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(13);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(12);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(11);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(10);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(9);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(8);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(7);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(6);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(5);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(4);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(3);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(2);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(1);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(0);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(15);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(14);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(13);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(12);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(11);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(10);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(9);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(8);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(7);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(6);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(5);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(4);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(3);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(2);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(1);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100100" |
                                   "100101" =>
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData37(0)
                                       & readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData21(0)
                                       & readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "100100" |
                                   "100101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2496 =>
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(15);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(14);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(13);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(12);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(11);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(10);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(9);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(8);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(7);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(6);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(5);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(4);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(3);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(2);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(1);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(0);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(15);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(14);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(13);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(12);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(11);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(10);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(9);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(8);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(7);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(6);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(5);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(4);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(3);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(2);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(1);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100100" |
                                   "100101" =>
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100110" =>
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData38(0)
                                       & readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData22(0)
                                       & readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "100100" |
                                   "100101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "100110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2560 =>
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "001";    
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(15);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(14);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(13);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(12);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(11);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(10);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(9);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(8);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(7);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(6);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(5);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(4);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(3);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(2);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(1);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(0);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(15);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(14);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(13);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(12);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(11);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(10);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(9);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(8);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(7);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(6);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(5);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(4);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(3);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(2);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(1);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(0);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData0_xhdl219 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData39(0)
                                       & readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData23(0)
                                       & readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData7(1 
                                       DOWNTO 0) & readData6(1 DOWNTO 0) 
                                       & readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0) & 
                                       readData0(1 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2624 =>
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "100";    
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(15);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(14);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(13);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(12);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(11);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(10);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(9);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(8);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(7);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(6);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(5);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(4);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(3);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(2);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(1);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(0);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(15);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(14);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(13);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(12);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(11);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(10);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(9);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(8);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(7);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(6);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(5);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(4);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(3);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(2);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(1);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(0);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" =>
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData40(0)
                                       & readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData24(0)
                                       & readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData8(1 
                                       DOWNTO 0) & readData7(1 DOWNTO 0) 
                                       & readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0);    
                              WHEN "101000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2688 =>
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(15);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(14);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(13);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(12);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(11);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(10);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(9);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(8);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(7);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(6);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(5);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(4);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(3);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(2);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(1);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(0);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(15);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(14);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(13);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(12);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(11);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(10);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(9);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(8);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(7);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(6);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(5);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(4);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(3);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(2);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(1);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(0);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" |
                                   "101001" =>
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData41(0)
                                       & readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData25(0)
                                       & readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData9(1 
                                       DOWNTO 0) & readData8(1 DOWNTO 0) 
                                       & readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0);    
                              WHEN "101000" |
                                   "101001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2752 =>
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(15);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(14);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(13);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(12);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(11);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(10);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(9);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(8);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(7);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(6);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(5);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(4);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(3);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(2);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(1);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(0);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(15);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(14);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(13);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(12);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(11);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(10);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(9);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(8);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(7);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(6);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(5);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(4);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(3);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(2);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(1);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(0);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" |
                                   "101001" =>
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101010" =>
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData42(0)
                                       & readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData26(0)
                                       & readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData10(1 
                                       DOWNTO 0) & readData9(1 DOWNTO 0) 
                                       & readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0);    
                              WHEN "101000" |
                                   "101001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "101010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2816 =>
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(15);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(14);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(13);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(12);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(11);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(10);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(9);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(8);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(7);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(6);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(5);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(4);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(3);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(2);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(1);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(0);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(15);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(14);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(13);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(12);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(11);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(10);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(9);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(8);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(7);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(6);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(5);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(4);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(3);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(2);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(1);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(0);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData43(0)
                                       & readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData27(0)
                                       & readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData11(1 
                                       DOWNTO 0) & readData10(1 DOWNTO 0)
                                       & readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0);    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2880 =>
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(15);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(14);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(13);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(12);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(11);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(10);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(9);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(8);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(7);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(6);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(5);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(4);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(3);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(2);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(1);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(0);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(15);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(14);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(13);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(12);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(11);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(10);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(9);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(8);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(7);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(6);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(5);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(4);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(3);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(2);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(1);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(0);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101100" =>
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData44(0)
                                       & readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData28(0)
                                       & readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData12(1 
                                       DOWNTO 0) & readData11(1 DOWNTO 0)
                                       & readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0);    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "101100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 2944 =>
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(15);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(14);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(13);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(12);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(11);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(10);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(9);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(8);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(7);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(6);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(5);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(4);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(3);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(2);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(1);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(0);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(15);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(14);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(13);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(12);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(11);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(10);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(9);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(8);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(7);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(6);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(5);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(4);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(3);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(2);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(1);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(0);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101100" |
                                   "101101" =>
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData45(0)
                                       & readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData29(0)
                                       & readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData13(1 
                                       DOWNTO 0) & readData12(1 DOWNTO 0)
                                       & readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0);    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "101100" |
                                   "101101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3008 =>
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "001";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(15);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(14);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(13);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(12);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(11);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(10);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(9);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(8);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(7);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(6);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(5);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(4);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(3);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(2);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(1);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(0);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(15);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(14);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(13);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(12);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(11);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(10);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(9);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(8);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(7);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(6);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(5);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(4);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(3);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(2);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(1);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(0);    
                           writeData14_xhdl233 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101100" |
                                   "101101" =>
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "101110" =>
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData46(0)
                                       & readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData30(0)
                                       & readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData14(1 
                                       DOWNTO 0) & readData13(1 DOWNTO 0)
                                       & readData12(1 DOWNTO 0) & 
                                       readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0);    
                              WHEN "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "101100" |
                                   "101101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "101110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3072 =>
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "000";    
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(9 DOWNTO 0);  
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(9 DOWNTO 0);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(15);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(14);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(13);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(12);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(11);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(10);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(9);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(8);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(7);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(6);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(5);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(4);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(3);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(2);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(1);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(0);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(15);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(14);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(13);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(12);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(11);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(10);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(9);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(8);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(7);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(6);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(5);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(4);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(3);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(2);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(1);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(0);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(15);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(14);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(13);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(12);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(11);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(10);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(9);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(8);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(7);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(6);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(5);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(4);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(3);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(2);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(1);    
                           writeData0_xhdl219 := "00000000000000000" & 
                           writeData(0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData47(0)
                                       & readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData31(0)
                                       & readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData15(0)
                                       & readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0) & readData1(0) & 
                                       readData0(0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3136 =>
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "100";    
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(15);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(14);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(13);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(12);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(11);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(10);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(9);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(8);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(7);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(6);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(5);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(4);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(3);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(2);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(1);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(0);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(15);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(14);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(13);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(12);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(11);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(10);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(9);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(8);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(7);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(6);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(5);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(4);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(3);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(2);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(1);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(0);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(15);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(14);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(13);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(12);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(11);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(10);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(9);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(8);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(7);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(6);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(5);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(4);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(3);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(2);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(1);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" =>
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData48(0)
                                       & readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData32(0)
                                       & readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData16(0)
                                       & readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0) & readData2(0) & 
                                       readData1(0);    
                              WHEN "110000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3200 =>
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(15);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(14);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(13);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(12);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(11);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(10);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(9);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(8);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(7);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(6);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(5);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(4);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(3);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(2);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(1);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(0);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(15);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(14);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(13);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(12);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(11);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(10);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(9);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(8);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(7);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(6);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(5);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(4);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(3);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(2);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(1);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(0);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(15);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(14);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(13);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(12);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(11);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(10);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(9);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(8);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(7);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(6);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(5);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(4);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(3);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(2);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(1);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" =>
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData49(0)
                                       & readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData33(0)
                                       & readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData17(0)
                                       & readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0);    
                              WHEN "110000" |
                                   "110001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3264 =>
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(15);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(14);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(13);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(12);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(11);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(10);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(9);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(8);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(7);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(6);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(5);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(4);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(3);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(2);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(1);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(0);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(15);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(14);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(13);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(12);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(11);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(10);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(9);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(8);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(7);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(6);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(5);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(4);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(3);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(2);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(1);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(0);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(15);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(14);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(13);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(12);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(11);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(10);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(9);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(8);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(7);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(6);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(5);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(4);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(3);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(2);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(1);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" =>
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110010" =>
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData50(0)
                                       & readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData34(0)
                                       & readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData18(0)
                                       & readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0);    
                              WHEN "110000" |
                                   "110001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "110010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3328 =>
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(15);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(14);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(13);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(12);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(11);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(10);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(9);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(8);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(7);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(6);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(5);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(4);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(3);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(2);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(1);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(0);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(15);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(14);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(13);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(12);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(11);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(10);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(9);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(8);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(7);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(6);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(5);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(4);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(3);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(2);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(1);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(0);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(15);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(14);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(13);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(12);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(11);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(10);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(9);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(8);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(7);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(6);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(5);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(4);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(3);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(2);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(1);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData51(0)
                                       & readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData35(0)
                                       & readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData19(0)
                                       & readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3392 =>
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(15);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(14);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(13);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(12);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(11);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(10);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(9);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(8);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(7);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(6);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(5);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(4);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(3);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(2);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(1);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(0);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(15);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(14);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(13);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(12);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(11);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(10);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(9);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(8);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(7);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(6);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(5);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(4);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(3);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(2);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(1);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(0);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(15);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(14);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(13);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(12);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(11);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(10);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(9);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(8);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(7);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(6);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(5);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(4);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(3);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(2);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(1);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110100" =>
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData52(0)
                                       & readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData36(0)
                                       & readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData20(0)
                                       & readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "110100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3456 =>
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(15);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(14);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(13);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(12);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(11);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(10);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(9);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(8);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(7);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(6);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(5);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(4);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(3);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(2);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(1);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(0);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(15);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(14);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(13);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(12);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(11);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(10);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(9);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(8);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(7);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(6);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(5);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(4);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(3);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(2);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(1);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(0);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(15);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(14);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(13);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(12);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(11);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(10);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(9);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(8);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(7);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(6);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(5);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(4);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(3);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(2);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(1);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110100" |
                                   "110101" =>
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData53(0)
                                       & readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData37(0)
                                       & readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData21(0)
                                       & readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "110100" |
                                   "110101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3520 =>
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(15);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(14);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(13);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(12);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(11);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(10);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(9);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(8);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(7);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(6);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(5);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(4);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(3);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(2);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(1);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(0);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(15);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(14);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(13);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(12);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(11);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(10);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(9);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(8);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(7);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(6);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(5);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(4);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(3);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(2);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(1);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(0);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(15);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(14);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(13);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(12);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(11);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(10);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(9);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(8);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(7);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(6);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(5);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(4);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(3);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(2);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(1);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110100" |
                                   "110101" =>
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110110" =>
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData54(0)
                                       & readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData38(0)
                                       & readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData22(0)
                                       & readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "110100" |
                                   "110101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "110110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3584 =>
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "001";    
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(15);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(14);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(13);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(12);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(11);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(10);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(9);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(8);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(7);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(6);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(5);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(4);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(3);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(2);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(1);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(0);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(15);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(14);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(13);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(12);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(11);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(10);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(9);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(8);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(7);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(6);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(5);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(4);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(3);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(2);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(1);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(0);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(15);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(14);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(13);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(12);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(11);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(10);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(9);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(8);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(7);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(6);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(5);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(4);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(3);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(2);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(1);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(0);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData0_xhdl219 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData55(0)
                                       & readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData39(0)
                                       & readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData23(0)
                                       & readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData7(1 
                                       DOWNTO 0) & readData6(1 DOWNTO 0) 
                                       & readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0) & 
                                       readData0(1 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3648 =>
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "100";    
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(15);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(14);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(13);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(12);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(11);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(10);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(9);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(8);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(7);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(6);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(5);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(4);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(3);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(2);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(1);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(0);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(15);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(14);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(13);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(12);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(11);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(10);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(9);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(8);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(7);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(6);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(5);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(4);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(3);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(2);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(1);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(0);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(15);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(14);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(13);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(12);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(11);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(10);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(9);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(8);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(7);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(6);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(5);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(4);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(3);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(2);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(1);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(0);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" =>
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData56(0)
                                       & readData55(0) & readData54(0) & 
                                       readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData40(0)
                                       & readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData24(0)
                                       & readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData8(1 
                                       DOWNTO 0) & readData7(1 DOWNTO 0) 
                                       & readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0);    
                              WHEN "111000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3712 =>
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(15);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(14);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(13);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(12);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(11);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(10);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(9);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(8);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(7);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(6);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(5);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(4);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(3);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(2);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(1);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(0);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(15);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(14);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(13);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(12);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(11);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(10);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(9);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(8);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(7);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(6);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(5);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(4);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(3);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(2);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(1);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(0);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(15);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(14);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(13);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(12);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(11);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(10);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(9);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(8);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(7);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(6);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(5);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(4);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(3);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(2);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(1);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(0);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" |
                                   "111001" =>
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData57(0)
                                       & readData56(0) & readData55(0) & 
                                       readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData41(0)
                                       & readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData25(0)
                                       & readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData9(1 
                                       DOWNTO 0) & readData8(1 DOWNTO 0) 
                                       & readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0);    
                              WHEN "111000" |
                                   "111001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3776 =>
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(15);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(14);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(13);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(12);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(11);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(10);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(9);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(8);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(7);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(6);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(5);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(4);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(3);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(2);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(1);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(0);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(15);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(14);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(13);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(12);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(11);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(10);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(9);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(8);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(7);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(6);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(5);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(4);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(3);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(2);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(1);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(0);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(15);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(14);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(13);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(12);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(11);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(10);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(9);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(8);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(7);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(6);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(5);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(4);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(3);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(2);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(1);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(0);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" |
                                   "111001" =>
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111010" =>
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData58(0)
                                       & readData57(0) & readData56(0) & 
                                       readData55(0) & readData54(0) & 
                                       readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData42(0)
                                       & readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData26(0)
                                       & readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData10(1 
                                       DOWNTO 0) & readData9(1 DOWNTO 0) 
                                       & readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0);    
                              WHEN "111000" |
                                   "111001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "111010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3840 =>
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(15);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(14);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(13);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(12);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(11);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(10);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(9);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(8);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(7);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(6);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(5);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(4);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(3);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(2);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(1);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(0);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(15);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(14);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(13);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(12);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(11);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(10);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(9);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(8);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(7);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(6);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(5);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(4);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(3);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(2);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(1);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(0);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(15);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(14);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(13);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(12);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(11);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(10);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(9);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(8);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(7);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(6);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(5);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(4);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(3);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(2);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(1);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(0);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData59(0)
                                       & readData58(0) & readData57(0) & 
                                       readData56(0) & readData55(0) & 
                                       readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData43(0)
                                       & readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData27(0)
                                       & readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData11(1 
                                       DOWNTO 0) & readData10(1 DOWNTO 0)
                                       & readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0);    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3904 =>
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(15);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(14);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(13);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(12);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(11);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(10);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(9);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(8);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(7);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(6);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(5);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(4);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(3);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(2);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(1);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(0);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(15);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(14);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(13);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(12);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(11);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(10);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(9);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(8);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(7);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(6);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(5);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(4);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(3);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(2);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(1);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(0);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(15);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(14);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(13);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(12);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(11);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(10);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(9);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(8);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(7);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(6);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(5);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(4);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(3);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(2);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(1);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(0);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111100" =>
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData60(0)
                                       & readData59(0) & readData58(0) & 
                                       readData57(0) & readData56(0) & 
                                       readData55(0) & readData54(0) & 
                                       readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData44(0)
                                       & readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData28(0)
                                       & readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData12(1 
                                       DOWNTO 0) & readData11(1 DOWNTO 0)
                                       & readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0) & 
                                       readData5(1 DOWNTO 0);    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "111100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 3968 =>
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(15);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(14);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(13);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(12);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(11);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(10);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(9);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(8);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(7);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(6);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(5);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(4);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(3);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(2);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(1);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(0);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(15);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(14);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(13);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(12);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(11);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(10);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(9);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(8);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(7);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(6);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(5);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(4);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(3);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(2);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(1);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(0);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(15);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(14);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(13);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(12);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(11);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(10);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(9);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(8);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(7);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(6);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(5);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(4);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(3);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(2);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(1);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(0);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111100" |
                                   "111101" =>
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData61(0)
                                       & readData60(0) & readData59(0) & 
                                       readData58(0) & readData57(0) & 
                                       readData56(0) & readData55(0) & 
                                       readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData45(0)
                                       & readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData29(0)
                                       & readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData13(1 
                                       DOWNTO 0) & readData12(1 DOWNTO 0)
                                       & readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0) & 
                                       readData6(1 DOWNTO 0);    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "111100" |
                                   "111101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4032 =>
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "001";    
                           width13_xhdl16 := "001";    
                           width12_xhdl15 := "001";    
                           width11_xhdl14 := "001";    
                           width10_xhdl13 := "001";    
                           width9_xhdl12 := "001";    
                           width8_xhdl11 := "001";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr13_xhdl304 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr12_xhdl303 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr11_xhdl302 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr10_xhdl301 := writeAddr(8 DOWNTO 0) 
                           & '0';    
                           writeAddr9_xhdl300 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr8_xhdl299 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr13_xhdl376 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr12_xhdl375 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr11_xhdl374 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr10_xhdl373 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr9_xhdl372 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr8_xhdl371 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(15);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(14);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(13);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(12);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(11);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(10);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(9);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(8);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(7);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(6);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(5);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(4);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(3);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(2);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(1);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(0);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(15);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(14);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(13);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(12);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(11);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(10);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(9);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(8);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(7);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(6);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(5);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(4);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(3);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(2);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(1);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(0);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(15);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(14);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(13);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(12);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(11);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(10);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(9);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(8);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(7);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(6);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(5);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(4);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(3);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(2);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(1);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(0);    
                           writeData14_xhdl233 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData13_xhdl232 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData12_xhdl231 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData11_xhdl230 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData10_xhdl229 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData9_xhdl228 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData8_xhdl227 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111100" |
                                   "111101" =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "111110" =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData62(0)
                                       & readData61(0) & readData60(0) & 
                                       readData59(0) & readData58(0) & 
                                       readData57(0) & readData56(0) & 
                                       readData55(0) & readData54(0) & 
                                       readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData46(0)
                                       & readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData30(0)
                                       & readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData14(1 
                                       DOWNTO 0) & readData13(1 DOWNTO 0)
                                       & readData12(1 DOWNTO 0) & 
                                       readData11(1 DOWNTO 0) & 
                                       readData10(1 DOWNTO 0) & 
                                       readData9(1 DOWNTO 0) & 
                                       readData8(1 DOWNTO 0) & 
                                       readData7(1 DOWNTO 0);    
                              WHEN "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "111100" |
                                   "111101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "111110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4096 =>
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "000";    
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(9 DOWNTO 0);  
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(9 DOWNTO 0);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(15);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(14);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(13);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(12);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(11);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(10);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(9);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(8);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(7);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(6);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(5);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(4);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(3);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(2);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(1);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(0);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(15);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(14);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(13);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(12);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(11);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(10);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(9);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(8);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(7);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(6);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(5);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(4);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(3);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(2);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(1);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(0);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(15);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(14);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(13);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(12);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(11);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(10);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(9);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(8);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(7);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(6);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(5);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(4);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(3);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(2);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(1);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(0);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(15);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(14);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(13);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(12);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(11);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(10);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(9);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(8);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(7);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(6);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(5);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(4);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(3);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(2);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(1);    
                           writeData0_xhdl219 := "00000000000000000" & 
                           writeData(0);    
                           CASE writeAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" |
                                   "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" |
                                   "111100" |
                                   "111101" |
                                   "111110" |
                                   "111111" =>
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(11 DOWNTO 6) IS
                              WHEN "000000" |
                                   "000001" |
                                   "000010" |
                                   "000011" |
                                   "000100" |
                                   "000101" |
                                   "000110" |
                                   "000111" |
                                   "001000" |
                                   "001001" |
                                   "001010" |
                                   "001011" |
                                   "001100" |
                                   "001101" |
                                   "001110" |
                                   "001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData63(0)
                                       & readData62(0) & readData61(0) & 
                                       readData60(0) & readData59(0) & 
                                       readData58(0) & readData57(0) & 
                                       readData56(0) & readData55(0) & 
                                       readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0);    
                              -- case: 6'b000000, 6'b000001, 6'b000010, 6'b000011, 6'b000100, 6'b000101,6'b000110, 6'b000111, 6'b001000, 6'b001001,...
                              
                              WHEN "010000" |
                                   "010001" |
                                   "010010" |
                                   "010011" |
                                   "010100" |
                                   "010101" |
                                   "010110" |
                                   "010111" |
                                   "011000" |
                                   "011001" |
                                   "011010" |
                                   "011011" |
                                   "011100" |
                                   "011101" |
                                   "011110" |
                                   "011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData47(0)
                                       & readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0);    
                              WHEN "100000" |
                                   "100001" |
                                   "100010" |
                                   "100011" |
                                   "100100" |
                                   "100101" |
                                   "100110" |
                                   "100111" |
                                   "101000" |
                                   "101001" |
                                   "101010" |
                                   "101011" |
                                   "101100" |
                                   "101101" |
                                   "101110" |
                                   "101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData31(0)
                                       & readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0);    
                              WHEN "110000" |
                                   "110001" |
                                   "110010" |
                                   "110011" |
                                   "110100" |
                                   "110101" |
                                   "110110" |
                                   "110111" |
                                   "111000" |
                                   "111001" |
                                   "111010" |
                                   "111011" |
                                   "111100" |
                                   "111101" |
                                   "111110" |
                                   "111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData15(0)
                                       & readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0) & readData1(0) & 
                                       readData0(0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4160 =>
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "000";    
                           width0_xhdl3 := "100";    
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(9 DOWNTO 0);  
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(9 DOWNTO 0);    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(15);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(14);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(13);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(12);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(11);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(10);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(9);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(8);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(7);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(6);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(5);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(4);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(3);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(2);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(1);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(0);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(15);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(14);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(13);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(12);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(11);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(10);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(9);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(8);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(7);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(6);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(5);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(4);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(3);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(2);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(1);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(0);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(15);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(14);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(13);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(12);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(11);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(10);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(9);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(8);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(7);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(6);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(5);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(4);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(3);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(2);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(1);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(0);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(15);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(14);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(13);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(12);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(11);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(10);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(9);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(8);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(7);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(6);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(5);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(4);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(3);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(2);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(1);    
                           writeData1_xhdl220 := "00000000000000000" & 
                           writeData(0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" =>
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData64(0)
                                       & readData63(0) & readData62(0) & 
                                       readData61(0) & readData60(0) & 
                                       readData59(0) & readData58(0) & 
                                       readData57(0) & readData56(0) & 
                                       readData55(0) & readData54(0) & 
                                       readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData48(0)
                                       & readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData32(0)
                                       & readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData16(0)
                                       & readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0) & readData2(0) & 
                                       readData1(0);    
                              WHEN "1000000" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4224 =>
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "000";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(9 DOWNTO 0);  
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(9 DOWNTO 0);    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(15);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(14);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(13);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(12);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(11);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(10);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(9);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(8);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(7);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(6);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(5);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(4);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(3);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(2);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(1);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(0);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(15);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(14);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(13);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(12);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(11);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(10);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(9);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(8);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(7);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(6);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(5);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(4);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(3);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(2);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(1);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(0);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(15);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(14);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(13);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(12);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(11);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(10);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(9);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(8);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(7);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(6);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(5);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(4);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(3);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(2);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(1);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(0);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(15);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(14);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(13);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(12);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(11);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(10);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(9);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(8);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(7);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(6);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(5);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(4);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(3);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(2);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(1);    
                           writeData2_xhdl221 := "00000000000000000" & 
                           writeData(0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" =>
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData65(0)
                                       & readData64(0) & readData63(0) & 
                                       readData62(0) & readData61(0) & 
                                       readData60(0) & readData59(0) & 
                                       readData58(0) & readData57(0) & 
                                       readData56(0) & readData55(0) & 
                                       readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData49(0)
                                       & readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData33(0)
                                       & readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData17(0)
                                       & readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0) & readData3(0) & 
                                       readData2(0);    
                              WHEN "1000000" |
                                   "1000001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4288 =>
                           width66_xhdl69 := "000";    
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "000";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr66_xhdl357 := writeAddr(9 DOWNTO 0); 
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(9 DOWNTO 0);  
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr66_xhdl429 := readAddr(9 DOWNTO 0);   
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(9 DOWNTO 0);    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData66_xhdl285 := "00000000000000000" & 
                           writeData(15);    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(14);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(13);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(12);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(11);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(10);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(9);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(8);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(7);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(6);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(5);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(4);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(3);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(2);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(1);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(0);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(15);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(14);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(13);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(12);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(11);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(10);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(9);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(8);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(7);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(6);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(5);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(4);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(3);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(2);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(1);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(0);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(15);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(14);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(13);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(12);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(11);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(10);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(9);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(8);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(7);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(6);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(5);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(4);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(3);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(2);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(1);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(0);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(15);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(14);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(13);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(12);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(11);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(10);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(9);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(8);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(7);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(6);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(5);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(4);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(3);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(2);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(1);    
                           writeData3_xhdl222 := "00000000000000000" & 
                           writeData(0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a66_xhdl141 := wen;    
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" =>
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000010" =>
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData66(0)
                                       & readData65(0) & readData64(0) & 
                                       readData63(0) & readData62(0) & 
                                       readData61(0) & readData60(0) & 
                                       readData59(0) & readData58(0) & 
                                       readData57(0) & readData56(0) & 
                                       readData55(0) & readData54(0) & 
                                       readData53(0) & readData52(0) & 
                                       readData51(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData50(0)
                                       & readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0) & readData36(0) & 
                                       readData35(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData34(0)
                                       & readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0) & readData20(0) & 
                                       readData19(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData18(0)
                                       & readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0) & readData4(0) & 
                                       readData3(0);    
                              WHEN "1000000" |
                                   "1000001" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "1000010" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4352 =>
                           width67_xhdl70 := "000";    
                           width66_xhdl69 := "000";    
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "000";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "010";    
                           writeAddr67_xhdl358 := writeAddr(9 DOWNTO 0); 
                           writeAddr66_xhdl357 := writeAddr(9 DOWNTO 0); 
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(9 DOWNTO 0);  
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr67_xhdl430 := readAddr(9 DOWNTO 0);   
                           readAddr66_xhdl429 := readAddr(9 DOWNTO 0);   
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(9 DOWNTO 0);    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           writeData67_xhdl286 := "00000000000000000" & 
                           writeData(15);    
                           writeData66_xhdl285 := "00000000000000000" & 
                           writeData(14);    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(13);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(12);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(11);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(10);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(9);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(8);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(7);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(6);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(5);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(4);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(3);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(2);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(1);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(0);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(15);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(14);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(13);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(12);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(11);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(10);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(9);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(8);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(7);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(6);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(5);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(4);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(3);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(2);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(1);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(0);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(15);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(14);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(13);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(12);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(11);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(10);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(9);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(8);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(7);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(6);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(5);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(4);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(3);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(2);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(1);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(0);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(15);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(14);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(13);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(12);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(11);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(10);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(9);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(8);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(7);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(6);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(5);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(4);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(3);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(2);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(1);    
                           writeData4_xhdl223 := "00000000000000000" & 
                           writeData(0);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData0_xhdl219 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a67_xhdl142 := wen;    
                                       wen_a66_xhdl141 := wen;    
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData67(0)
                                       & readData66(0) & readData65(0) & 
                                       readData64(0) & readData63(0) & 
                                       readData62(0) & readData61(0) & 
                                       readData60(0) & readData59(0) & 
                                       readData58(0) & readData57(0) & 
                                       readData56(0) & readData55(0) & 
                                       readData54(0) & readData53(0) & 
                                       readData52(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData51(0)
                                       & readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0) & readData37(0) & 
                                       readData36(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData35(0)
                                       & readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0) & readData21(0) & 
                                       readData20(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData19(0)
                                       & readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0) & readData5(0) & 
                                       readData4(0);    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData3(3 
                                       DOWNTO 0) & readData2(3 DOWNTO 0) 
                                       & readData1(3 DOWNTO 0) & 
                                       readData0(3 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4416 =>
                           width68_xhdl71 := "000";    
                           width67_xhdl70 := "000";    
                           width66_xhdl69 := "000";    
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "000";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "010";    
                           width0_xhdl3 := "100";    
                           writeAddr68_xhdl359 := writeAddr(9 DOWNTO 0); 
                           writeAddr67_xhdl358 := writeAddr(9 DOWNTO 0); 
                           writeAddr66_xhdl357 := writeAddr(9 DOWNTO 0); 
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(9 DOWNTO 0);  
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr68_xhdl431 := readAddr(9 DOWNTO 0);   
                           readAddr67_xhdl430 := readAddr(9 DOWNTO 0);   
                           readAddr66_xhdl429 := readAddr(9 DOWNTO 0);   
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(9 DOWNTO 0);    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData68_xhdl287 := "00000000000000000" & 
                           writeData(15);    
                           writeData67_xhdl286 := "00000000000000000" & 
                           writeData(14);    
                           writeData66_xhdl285 := "00000000000000000" & 
                           writeData(13);    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(12);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(11);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(10);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(9);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(8);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(7);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(6);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(5);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(4);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(3);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(2);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(1);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(0);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(15);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(14);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(13);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(12);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(11);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(10);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(9);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(8);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(7);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(6);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(5);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(4);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(3);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(2);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(1);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(0);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(15);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(14);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(13);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(12);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(11);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(10);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(9);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(8);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(7);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(6);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(5);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(4);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(3);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(2);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(1);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(0);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(15);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(14);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(13);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(12);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(11);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(10);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(9);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(8);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(7);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(6);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(5);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(4);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(3);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(2);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(1);    
                           writeData5_xhdl224 := "00000000000000000" & 
                           writeData(0);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData1_xhdl220 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a68_xhdl143 := wen;    
                                       wen_a67_xhdl142 := wen;    
                                       wen_a66_xhdl141 := wen;    
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000100" =>
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData68(0)
                                       & readData67(0) & readData66(0) & 
                                       readData65(0) & readData64(0) & 
                                       readData63(0) & readData62(0) & 
                                       readData61(0) & readData60(0) & 
                                       readData59(0) & readData58(0) & 
                                       readData57(0) & readData56(0) & 
                                       readData55(0) & readData54(0) & 
                                       readData53(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData52(0)
                                       & readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0) & readData38(0) & 
                                       readData37(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData36(0)
                                       & readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0) & readData22(0) & 
                                       readData21(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData20(0)
                                       & readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0) & readData6(0) & 
                                       readData5(0);    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData4(3 
                                       DOWNTO 0) & readData3(3 DOWNTO 0) 
                                       & readData2(3 DOWNTO 0) & 
                                       readData1(3 DOWNTO 0);    
                              WHEN "1000100" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4480 =>
                           width69_xhdl72 := "000";    
                           width68_xhdl71 := "000";    
                           width67_xhdl70 := "000";    
                           width66_xhdl69 := "000";    
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "000";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "010";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "011";    
                           writeAddr69_xhdl360 := writeAddr(9 DOWNTO 0); 
                           writeAddr68_xhdl359 := writeAddr(9 DOWNTO 0); 
                           writeAddr67_xhdl358 := writeAddr(9 DOWNTO 0); 
                           writeAddr66_xhdl357 := writeAddr(9 DOWNTO 0); 
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(9 DOWNTO 0);  
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr69_xhdl432 := readAddr(9 DOWNTO 0);   
                           readAddr68_xhdl431 := readAddr(9 DOWNTO 0);   
                           readAddr67_xhdl430 := readAddr(9 DOWNTO 0);   
                           readAddr66_xhdl429 := readAddr(9 DOWNTO 0);   
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(9 DOWNTO 0);    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           writeData69_xhdl288 := "00000000000000000" & 
                           writeData(15);    
                           writeData68_xhdl287 := "00000000000000000" & 
                           writeData(14);    
                           writeData67_xhdl286 := "00000000000000000" & 
                           writeData(13);    
                           writeData66_xhdl285 := "00000000000000000" & 
                           writeData(12);    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(11);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(10);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(9);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(8);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(7);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(6);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(5);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(4);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(3);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(2);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(1);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(0);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(15);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(14);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(13);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(12);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(11);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(10);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(9);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(8);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(7);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(6);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(5);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(4);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(3);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(2);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(1);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(0);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(15);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(14);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(13);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(12);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(11);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(10);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(9);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(8);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(7);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(6);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(5);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(4);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(3);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(2);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(1);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(0);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(15);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(14);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(13);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(12);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(11);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(10);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(9);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(8);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(7);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(6);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(5);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(4);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(3);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(2);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(1);    
                           writeData6_xhdl225 := "00000000000000000" & 
                           writeData(0);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData2_xhdl221 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData0_xhdl219 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a69_xhdl144 := wen;    
                                       wen_a68_xhdl143 := wen;    
                                       wen_a67_xhdl142 := wen;    
                                       wen_a66_xhdl141 := wen;    
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000100" |
                                   "1000101" =>
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData69(0)
                                       & readData68(0) & readData67(0) & 
                                       readData66(0) & readData65(0) & 
                                       readData64(0) & readData63(0) & 
                                       readData62(0) & readData61(0) & 
                                       readData60(0) & readData59(0) & 
                                       readData58(0) & readData57(0) & 
                                       readData56(0) & readData55(0) & 
                                       readData54(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData53(0)
                                       & readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0) & readData39(0) & 
                                       readData38(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData37(0)
                                       & readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0) & readData23(0) & 
                                       readData22(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData21(0)
                                       & readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0) & readData7(0) & 
                                       readData6(0);    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData5(3 
                                       DOWNTO 0) & readData4(3 DOWNTO 0) 
                                       & readData3(3 DOWNTO 0) & 
                                       readData2(3 DOWNTO 0);    
                              WHEN "1000100" |
                                   "1000101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData1(7 
                                       DOWNTO 0) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4544 =>
                           width70_xhdl73 := "000";    
                           width69_xhdl72 := "000";    
                           width68_xhdl71 := "000";    
                           width67_xhdl70 := "000";    
                           width66_xhdl69 := "000";    
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "000";    
                           width6_xhdl9 := "010";    
                           width5_xhdl8 := "010";    
                           width4_xhdl7 := "010";    
                           width3_xhdl6 := "010";    
                           width2_xhdl5 := "011";    
                           width1_xhdl4 := "011";    
                           width0_xhdl3 := "100";    
                           writeAddr70_xhdl361 := writeAddr(9 DOWNTO 0); 
                           writeAddr69_xhdl360 := writeAddr(9 DOWNTO 0); 
                           writeAddr68_xhdl359 := writeAddr(9 DOWNTO 0); 
                           writeAddr67_xhdl358 := writeAddr(9 DOWNTO 0); 
                           writeAddr66_xhdl357 := writeAddr(9 DOWNTO 0); 
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(9 DOWNTO 0);  
                           writeAddr6_xhdl297 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr5_xhdl296 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr4_xhdl295 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr3_xhdl294 := writeAddr(7 DOWNTO 0) & 
                           "00";    
                           writeAddr2_xhdl293 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr1_xhdl292 := writeAddr(6 DOWNTO 0) & 
                           "000";    
                           writeAddr0_xhdl291 := writeAddr(5 DOWNTO 0) & 
                           "0000";    
                           readAddr70_xhdl433 := readAddr(9 DOWNTO 0);   
                           readAddr69_xhdl432 := readAddr(9 DOWNTO 0);   
                           readAddr68_xhdl431 := readAddr(9 DOWNTO 0);   
                           readAddr67_xhdl430 := readAddr(9 DOWNTO 0);   
                           readAddr66_xhdl429 := readAddr(9 DOWNTO 0);   
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(9 DOWNTO 0);    
                           readAddr6_xhdl369 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr5_xhdl368 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr4_xhdl367 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr3_xhdl366 := readAddr(7 DOWNTO 0) & 
                           "00";    
                           readAddr2_xhdl365 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr1_xhdl364 := readAddr(6 DOWNTO 0) & 
                           "000";    
                           readAddr0_xhdl363 := readAddr(5 DOWNTO 0) & 
                           "0000";    
                           writeData70_xhdl289 := "00000000000000000" & 
                           writeData(15);    
                           writeData69_xhdl288 := "00000000000000000" & 
                           writeData(14);    
                           writeData68_xhdl287 := "00000000000000000" & 
                           writeData(13);    
                           writeData67_xhdl286 := "00000000000000000" & 
                           writeData(12);    
                           writeData66_xhdl285 := "00000000000000000" & 
                           writeData(11);    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(10);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(9);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(8);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(7);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(6);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(5);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(4);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(3);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(2);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(1);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(0);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(15);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(14);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(13);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(12);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(11);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(10);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(9);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(8);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(7);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(6);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(5);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(4);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(3);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(2);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(1);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(0);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(15);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(14);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(13);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(12);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(11);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(10);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(9);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(8);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(7);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(6);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(5);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(4);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(3);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(2);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(1);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(0);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(15);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(14);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(13);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(12);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(11);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(10);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(9);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(8);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(7);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(6);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(5);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(4);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(3);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(2);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(1);    
                           writeData7_xhdl226 := "00000000000000000" & 
                           writeData(0);    
                           writeData6_xhdl225 := "00000000000000" & 
                           writeData(15 DOWNTO 12);    
                           writeData5_xhdl224 := "00000000000000" & 
                           writeData(11 DOWNTO 8);    
                           writeData4_xhdl223 := "00000000000000" & 
                           writeData(7 DOWNTO 4);    
                           writeData3_xhdl222 := "00000000000000" & 
                           writeData(3 DOWNTO 0);    
                           writeData2_xhdl221 := "0000000000" & 
                           writeData(15 DOWNTO 8);    
                           writeData1_xhdl220 := "0000000000" & 
                           writeData(7 DOWNTO 0);    
                           writeData0_xhdl219 := '0' & writeData(15 
                           DOWNTO 8) & '0' & writeData(7 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a70_xhdl145 := wen;    
                                       wen_a69_xhdl144 := wen;    
                                       wen_a68_xhdl143 := wen;    
                                       wen_a67_xhdl142 := wen;    
                                       wen_a66_xhdl141 := wen;    
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000100" |
                                   "1000101" =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000110" =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData70(0)
                                       & readData69(0) & readData68(0) & 
                                       readData67(0) & readData66(0) & 
                                       readData65(0) & readData64(0) & 
                                       readData63(0) & readData62(0) & 
                                       readData61(0) & readData60(0) & 
                                       readData59(0) & readData58(0) & 
                                       readData57(0) & readData56(0) & 
                                       readData55(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData54(0)
                                       & readData53(0) & readData52(0) & 
                                       readData51(0) & readData50(0) & 
                                       readData49(0) & readData48(0) & 
                                       readData47(0) & readData46(0) & 
                                       readData45(0) & readData44(0) & 
                                       readData43(0) & readData42(0) & 
                                       readData41(0) & readData40(0) & 
                                       readData39(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData38(0)
                                       & readData37(0) & readData36(0) & 
                                       readData35(0) & readData34(0) & 
                                       readData33(0) & readData32(0) & 
                                       readData31(0) & readData30(0) & 
                                       readData29(0) & readData28(0) & 
                                       readData27(0) & readData26(0) & 
                                       readData25(0) & readData24(0) & 
                                       readData23(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData22(0)
                                       & readData21(0) & readData20(0) & 
                                       readData19(0) & readData18(0) & 
                                       readData17(0) & readData16(0) & 
                                       readData15(0) & readData14(0) & 
                                       readData13(0) & readData12(0) & 
                                       readData11(0) & readData10(0) & 
                                       readData9(0) & readData8(0) & 
                                       readData7(0);    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData6(3 
                                       DOWNTO 0) & readData5(3 DOWNTO 0) 
                                       & readData4(3 DOWNTO 0) & 
                                       readData3(3 DOWNTO 0);    
                              WHEN "1000100" |
                                   "1000101" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData2(7 
                                       DOWNTO 0) & readData1(7 DOWNTO 0)
                                       ;    
                              WHEN "1000110" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData0(16 
                                       DOWNTO 9) & readData0(7 DOWNTO 0)
                                       ;    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN 4608 =>
                           width71_xhdl74 := "000";    
                           width70_xhdl73 := "000";    
                           width69_xhdl72 := "000";    
                           width68_xhdl71 := "000";    
                           width67_xhdl70 := "000";    
                           width66_xhdl69 := "000";    
                           width65_xhdl68 := "000";    
                           width64_xhdl67 := "000";    
                           width63_xhdl66 := "000";    
                           width62_xhdl65 := "000";    
                           width61_xhdl64 := "000";    
                           width60_xhdl63 := "000";    
                           width59_xhdl62 := "000";    
                           width58_xhdl61 := "000";    
                           width57_xhdl60 := "000";    
                           width56_xhdl59 := "000";    
                           width55_xhdl58 := "000";    
                           width54_xhdl57 := "000";    
                           width53_xhdl56 := "000";    
                           width52_xhdl55 := "000";    
                           width51_xhdl54 := "000";    
                           width50_xhdl53 := "000";    
                           width49_xhdl52 := "000";    
                           width48_xhdl51 := "000";    
                           width47_xhdl50 := "000";    
                           width46_xhdl49 := "000";    
                           width45_xhdl48 := "000";    
                           width44_xhdl47 := "000";    
                           width43_xhdl46 := "000";    
                           width42_xhdl45 := "000";    
                           width41_xhdl44 := "000";    
                           width40_xhdl43 := "000";    
                           width39_xhdl42 := "000";    
                           width38_xhdl41 := "000";    
                           width37_xhdl40 := "000";    
                           width36_xhdl39 := "000";    
                           width35_xhdl38 := "000";    
                           width34_xhdl37 := "000";    
                           width33_xhdl36 := "000";    
                           width32_xhdl35 := "000";    
                           width31_xhdl34 := "000";    
                           width30_xhdl33 := "000";    
                           width29_xhdl32 := "000";    
                           width28_xhdl31 := "000";    
                           width27_xhdl30 := "000";    
                           width26_xhdl29 := "000";    
                           width25_xhdl28 := "000";    
                           width24_xhdl27 := "000";    
                           width23_xhdl26 := "000";    
                           width22_xhdl25 := "000";    
                           width21_xhdl24 := "000";    
                           width20_xhdl23 := "000";    
                           width19_xhdl22 := "000";    
                           width18_xhdl21 := "000";    
                           width17_xhdl20 := "000";    
                           width16_xhdl19 := "000";    
                           width15_xhdl18 := "000";    
                           width14_xhdl17 := "000";    
                           width13_xhdl16 := "000";    
                           width12_xhdl15 := "000";    
                           width11_xhdl14 := "000";    
                           width10_xhdl13 := "000";    
                           width9_xhdl12 := "000";    
                           width8_xhdl11 := "000";    
                           width7_xhdl10 := "001";    
                           width6_xhdl9 := "001";    
                           width5_xhdl8 := "001";    
                           width4_xhdl7 := "001";    
                           width3_xhdl6 := "001";    
                           width2_xhdl5 := "001";    
                           width1_xhdl4 := "001";    
                           width0_xhdl3 := "001";    
                           writeAddr71_xhdl362 := writeAddr(9 DOWNTO 0); 
                           writeAddr70_xhdl361 := writeAddr(9 DOWNTO 0); 
                           writeAddr69_xhdl360 := writeAddr(9 DOWNTO 0); 
                           writeAddr68_xhdl359 := writeAddr(9 DOWNTO 0); 
                           writeAddr67_xhdl358 := writeAddr(9 DOWNTO 0); 
                           writeAddr66_xhdl357 := writeAddr(9 DOWNTO 0); 
                           writeAddr65_xhdl356 := writeAddr(9 DOWNTO 0); 
                           writeAddr64_xhdl355 := writeAddr(9 DOWNTO 0); 
                           writeAddr63_xhdl354 := writeAddr(9 DOWNTO 0); 
                           writeAddr62_xhdl353 := writeAddr(9 DOWNTO 0); 
                           writeAddr61_xhdl352 := writeAddr(9 DOWNTO 0); 
                           writeAddr60_xhdl351 := writeAddr(9 DOWNTO 0); 
                           writeAddr59_xhdl350 := writeAddr(9 DOWNTO 0); 
                           writeAddr58_xhdl349 := writeAddr(9 DOWNTO 0); 
                           writeAddr57_xhdl348 := writeAddr(9 DOWNTO 0); 
                           writeAddr56_xhdl347 := writeAddr(9 DOWNTO 0); 
                           writeAddr55_xhdl346 := writeAddr(9 DOWNTO 0); 
                           writeAddr54_xhdl345 := writeAddr(9 DOWNTO 0); 
                           writeAddr53_xhdl344 := writeAddr(9 DOWNTO 0); 
                           writeAddr52_xhdl343 := writeAddr(9 DOWNTO 0); 
                           writeAddr51_xhdl342 := writeAddr(9 DOWNTO 0); 
                           writeAddr50_xhdl341 := writeAddr(9 DOWNTO 0); 
                           writeAddr49_xhdl340 := writeAddr(9 DOWNTO 0); 
                           writeAddr48_xhdl339 := writeAddr(9 DOWNTO 0); 
                           writeAddr47_xhdl338 := writeAddr(9 DOWNTO 0); 
                           writeAddr46_xhdl337 := writeAddr(9 DOWNTO 0); 
                           writeAddr45_xhdl336 := writeAddr(9 DOWNTO 0); 
                           writeAddr44_xhdl335 := writeAddr(9 DOWNTO 0); 
                           writeAddr43_xhdl334 := writeAddr(9 DOWNTO 0); 
                           writeAddr42_xhdl333 := writeAddr(9 DOWNTO 0); 
                           writeAddr41_xhdl332 := writeAddr(9 DOWNTO 0); 
                           writeAddr40_xhdl331 := writeAddr(9 DOWNTO 0); 
                           writeAddr39_xhdl330 := writeAddr(9 DOWNTO 0); 
                           writeAddr38_xhdl329 := writeAddr(9 DOWNTO 0); 
                           writeAddr37_xhdl328 := writeAddr(9 DOWNTO 0); 
                           writeAddr36_xhdl327 := writeAddr(9 DOWNTO 0); 
                           writeAddr35_xhdl326 := writeAddr(9 DOWNTO 0); 
                           writeAddr34_xhdl325 := writeAddr(9 DOWNTO 0); 
                           writeAddr33_xhdl324 := writeAddr(9 DOWNTO 0); 
                           writeAddr32_xhdl323 := writeAddr(9 DOWNTO 0); 
                           writeAddr31_xhdl322 := writeAddr(9 DOWNTO 0); 
                           writeAddr30_xhdl321 := writeAddr(9 DOWNTO 0); 
                           writeAddr29_xhdl320 := writeAddr(9 DOWNTO 0); 
                           writeAddr28_xhdl319 := writeAddr(9 DOWNTO 0); 
                           writeAddr27_xhdl318 := writeAddr(9 DOWNTO 0); 
                           writeAddr26_xhdl317 := writeAddr(9 DOWNTO 0); 
                           writeAddr25_xhdl316 := writeAddr(9 DOWNTO 0); 
                           writeAddr24_xhdl315 := writeAddr(9 DOWNTO 0); 
                           writeAddr23_xhdl314 := writeAddr(9 DOWNTO 0); 
                           writeAddr22_xhdl313 := writeAddr(9 DOWNTO 0); 
                           writeAddr21_xhdl312 := writeAddr(9 DOWNTO 0); 
                           writeAddr20_xhdl311 := writeAddr(9 DOWNTO 0); 
                           writeAddr19_xhdl310 := writeAddr(9 DOWNTO 0); 
                           writeAddr18_xhdl309 := writeAddr(9 DOWNTO 0); 
                           writeAddr17_xhdl308 := writeAddr(9 DOWNTO 0); 
                           writeAddr16_xhdl307 := writeAddr(9 DOWNTO 0); 
                           writeAddr15_xhdl306 := writeAddr(9 DOWNTO 0); 
                           writeAddr14_xhdl305 := writeAddr(9 DOWNTO 0); 
                           writeAddr13_xhdl304 := writeAddr(9 DOWNTO 0); 
                           writeAddr12_xhdl303 := writeAddr(9 DOWNTO 0); 
                           writeAddr11_xhdl302 := writeAddr(9 DOWNTO 0); 
                           writeAddr10_xhdl301 := writeAddr(9 DOWNTO 0); 
                           writeAddr9_xhdl300 := writeAddr(9 DOWNTO 0);  
                           writeAddr8_xhdl299 := writeAddr(9 DOWNTO 0);  
                           writeAddr7_xhdl298 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr6_xhdl297 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr5_xhdl296 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr4_xhdl295 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr3_xhdl294 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr2_xhdl293 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr1_xhdl292 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           writeAddr0_xhdl291 := writeAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr71_xhdl434 := readAddr(9 DOWNTO 0);   
                           readAddr70_xhdl433 := readAddr(9 DOWNTO 0);   
                           readAddr69_xhdl432 := readAddr(9 DOWNTO 0);   
                           readAddr68_xhdl431 := readAddr(9 DOWNTO 0);   
                           readAddr67_xhdl430 := readAddr(9 DOWNTO 0);   
                           readAddr66_xhdl429 := readAddr(9 DOWNTO 0);   
                           readAddr65_xhdl428 := readAddr(9 DOWNTO 0);   
                           readAddr64_xhdl427 := readAddr(9 DOWNTO 0);   
                           readAddr63_xhdl426 := readAddr(9 DOWNTO 0);   
                           readAddr62_xhdl425 := readAddr(9 DOWNTO 0);   
                           readAddr61_xhdl424 := readAddr(9 DOWNTO 0);   
                           readAddr60_xhdl423 := readAddr(9 DOWNTO 0);   
                           readAddr59_xhdl422 := readAddr(9 DOWNTO 0);   
                           readAddr58_xhdl421 := readAddr(9 DOWNTO 0);   
                           readAddr57_xhdl420 := readAddr(9 DOWNTO 0);   
                           readAddr56_xhdl419 := readAddr(9 DOWNTO 0);   
                           readAddr55_xhdl418 := readAddr(9 DOWNTO 0);   
                           readAddr54_xhdl417 := readAddr(9 DOWNTO 0);   
                           readAddr53_xhdl416 := readAddr(9 DOWNTO 0);   
                           readAddr52_xhdl415 := readAddr(9 DOWNTO 0);   
                           readAddr51_xhdl414 := readAddr(9 DOWNTO 0);   
                           readAddr50_xhdl413 := readAddr(9 DOWNTO 0);   
                           readAddr49_xhdl412 := readAddr(9 DOWNTO 0);   
                           readAddr48_xhdl411 := readAddr(9 DOWNTO 0);   
                           readAddr47_xhdl410 := readAddr(9 DOWNTO 0);   
                           readAddr46_xhdl409 := readAddr(9 DOWNTO 0);   
                           readAddr45_xhdl408 := readAddr(9 DOWNTO 0);   
                           readAddr44_xhdl407 := readAddr(9 DOWNTO 0);   
                           readAddr43_xhdl406 := readAddr(9 DOWNTO 0);   
                           readAddr42_xhdl405 := readAddr(9 DOWNTO 0);   
                           readAddr41_xhdl404 := readAddr(9 DOWNTO 0);   
                           readAddr40_xhdl403 := readAddr(9 DOWNTO 0);   
                           readAddr39_xhdl402 := readAddr(9 DOWNTO 0);   
                           readAddr38_xhdl401 := readAddr(9 DOWNTO 0);   
                           readAddr37_xhdl400 := readAddr(9 DOWNTO 0);   
                           readAddr36_xhdl399 := readAddr(9 DOWNTO 0);   
                           readAddr35_xhdl398 := readAddr(9 DOWNTO 0);   
                           readAddr34_xhdl397 := readAddr(9 DOWNTO 0);   
                           readAddr33_xhdl396 := readAddr(9 DOWNTO 0);   
                           readAddr32_xhdl395 := readAddr(9 DOWNTO 0);   
                           readAddr31_xhdl394 := readAddr(9 DOWNTO 0);   
                           readAddr30_xhdl393 := readAddr(9 DOWNTO 0);   
                           readAddr29_xhdl392 := readAddr(9 DOWNTO 0);   
                           readAddr28_xhdl391 := readAddr(9 DOWNTO 0);   
                           readAddr27_xhdl390 := readAddr(9 DOWNTO 0);   
                           readAddr26_xhdl389 := readAddr(9 DOWNTO 0);   
                           readAddr25_xhdl388 := readAddr(9 DOWNTO 0);   
                           readAddr24_xhdl387 := readAddr(9 DOWNTO 0);   
                           readAddr23_xhdl386 := readAddr(9 DOWNTO 0);   
                           readAddr22_xhdl385 := readAddr(9 DOWNTO 0);   
                           readAddr21_xhdl384 := readAddr(9 DOWNTO 0);   
                           readAddr20_xhdl383 := readAddr(9 DOWNTO 0);   
                           readAddr19_xhdl382 := readAddr(9 DOWNTO 0);   
                           readAddr18_xhdl381 := readAddr(9 DOWNTO 0);   
                           readAddr17_xhdl380 := readAddr(9 DOWNTO 0);   
                           readAddr16_xhdl379 := readAddr(9 DOWNTO 0);   
                           readAddr15_xhdl378 := readAddr(9 DOWNTO 0);   
                           readAddr14_xhdl377 := readAddr(9 DOWNTO 0);   
                           readAddr13_xhdl376 := readAddr(9 DOWNTO 0);   
                           readAddr12_xhdl375 := readAddr(9 DOWNTO 0);   
                           readAddr11_xhdl374 := readAddr(9 DOWNTO 0);   
                           readAddr10_xhdl373 := readAddr(9 DOWNTO 0);   
                           readAddr9_xhdl372 := readAddr(9 DOWNTO 0);    
                           readAddr8_xhdl371 := readAddr(9 DOWNTO 0);    
                           readAddr7_xhdl370 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr6_xhdl369 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr5_xhdl368 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr4_xhdl367 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr3_xhdl366 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr2_xhdl365 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr1_xhdl364 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           readAddr0_xhdl363 := readAddr(8 DOWNTO 0) & 
                           '0';    
                           writeData71_xhdl290 := "00000000000000000" & 
                           writeData(15);    
                           writeData70_xhdl289 := "00000000000000000" & 
                           writeData(14);    
                           writeData69_xhdl288 := "00000000000000000" & 
                           writeData(13);    
                           writeData68_xhdl287 := "00000000000000000" & 
                           writeData(12);    
                           writeData67_xhdl286 := "00000000000000000" & 
                           writeData(11);    
                           writeData66_xhdl285 := "00000000000000000" & 
                           writeData(10);    
                           writeData65_xhdl284 := "00000000000000000" & 
                           writeData(9);    
                           writeData64_xhdl283 := "00000000000000000" & 
                           writeData(8);    
                           writeData63_xhdl282 := "00000000000000000" & 
                           writeData(7);    
                           writeData62_xhdl281 := "00000000000000000" & 
                           writeData(6);    
                           writeData61_xhdl280 := "00000000000000000" & 
                           writeData(5);    
                           writeData60_xhdl279 := "00000000000000000" & 
                           writeData(4);    
                           writeData59_xhdl278 := "00000000000000000" & 
                           writeData(3);    
                           writeData58_xhdl277 := "00000000000000000" & 
                           writeData(2);    
                           writeData57_xhdl276 := "00000000000000000" & 
                           writeData(1);    
                           writeData56_xhdl275 := "00000000000000000" & 
                           writeData(0);    
                           writeData55_xhdl274 := "00000000000000000" & 
                           writeData(15);    
                           writeData54_xhdl273 := "00000000000000000" & 
                           writeData(14);    
                           writeData53_xhdl272 := "00000000000000000" & 
                           writeData(13);    
                           writeData52_xhdl271 := "00000000000000000" & 
                           writeData(12);    
                           writeData51_xhdl270 := "00000000000000000" & 
                           writeData(11);    
                           writeData50_xhdl269 := "00000000000000000" & 
                           writeData(10);    
                           writeData49_xhdl268 := "00000000000000000" & 
                           writeData(9);    
                           writeData48_xhdl267 := "00000000000000000" & 
                           writeData(8);    
                           writeData47_xhdl266 := "00000000000000000" & 
                           writeData(7);    
                           writeData46_xhdl265 := "00000000000000000" & 
                           writeData(6);    
                           writeData45_xhdl264 := "00000000000000000" & 
                           writeData(5);    
                           writeData44_xhdl263 := "00000000000000000" & 
                           writeData(4);    
                           writeData43_xhdl262 := "00000000000000000" & 
                           writeData(3);    
                           writeData42_xhdl261 := "00000000000000000" & 
                           writeData(2);    
                           writeData41_xhdl260 := "00000000000000000" & 
                           writeData(1);    
                           writeData40_xhdl259 := "00000000000000000" & 
                           writeData(0);    
                           writeData39_xhdl258 := "00000000000000000" & 
                           writeData(15);    
                           writeData38_xhdl257 := "00000000000000000" & 
                           writeData(14);    
                           writeData37_xhdl256 := "00000000000000000" & 
                           writeData(13);    
                           writeData36_xhdl255 := "00000000000000000" & 
                           writeData(12);    
                           writeData35_xhdl254 := "00000000000000000" & 
                           writeData(11);    
                           writeData34_xhdl253 := "00000000000000000" & 
                           writeData(10);    
                           writeData33_xhdl252 := "00000000000000000" & 
                           writeData(9);    
                           writeData32_xhdl251 := "00000000000000000" & 
                           writeData(8);    
                           writeData31_xhdl250 := "00000000000000000" & 
                           writeData(7);    
                           writeData30_xhdl249 := "00000000000000000" & 
                           writeData(6);    
                           writeData29_xhdl248 := "00000000000000000" & 
                           writeData(5);    
                           writeData28_xhdl247 := "00000000000000000" & 
                           writeData(4);    
                           writeData27_xhdl246 := "00000000000000000" & 
                           writeData(3);    
                           writeData26_xhdl245 := "00000000000000000" & 
                           writeData(2);    
                           writeData25_xhdl244 := "00000000000000000" & 
                           writeData(1);    
                           writeData24_xhdl243 := "00000000000000000" & 
                           writeData(0);    
                           writeData23_xhdl242 := "00000000000000000" & 
                           writeData(15);    
                           writeData22_xhdl241 := "00000000000000000" & 
                           writeData(14);    
                           writeData21_xhdl240 := "00000000000000000" & 
                           writeData(13);    
                           writeData20_xhdl239 := "00000000000000000" & 
                           writeData(12);    
                           writeData19_xhdl238 := "00000000000000000" & 
                           writeData(11);    
                           writeData18_xhdl237 := "00000000000000000" & 
                           writeData(10);    
                           writeData17_xhdl236 := "00000000000000000" & 
                           writeData(9);    
                           writeData16_xhdl235 := "00000000000000000" & 
                           writeData(8);    
                           writeData15_xhdl234 := "00000000000000000" & 
                           writeData(7);    
                           writeData14_xhdl233 := "00000000000000000" & 
                           writeData(6);    
                           writeData13_xhdl232 := "00000000000000000" & 
                           writeData(5);    
                           writeData12_xhdl231 := "00000000000000000" & 
                           writeData(4);    
                           writeData11_xhdl230 := "00000000000000000" & 
                           writeData(3);    
                           writeData10_xhdl229 := "00000000000000000" & 
                           writeData(2);    
                           writeData9_xhdl228 := "00000000000000000" & 
                           writeData(1);    
                           writeData8_xhdl227 := "00000000000000000" & 
                           writeData(0);    
                           writeData7_xhdl226 := "0000000000000000" & 
                           writeData(15 DOWNTO 14);    
                           writeData6_xhdl225 := "0000000000000000" & 
                           writeData(13 DOWNTO 12);    
                           writeData5_xhdl224 := "0000000000000000" & 
                           writeData(11 DOWNTO 10);    
                           writeData4_xhdl223 := "0000000000000000" & 
                           writeData(9 DOWNTO 8);    
                           writeData3_xhdl222 := "0000000000000000" & 
                           writeData(7 DOWNTO 6);    
                           writeData2_xhdl221 := "0000000000000000" & 
                           writeData(5 DOWNTO 4);    
                           writeData1_xhdl220 := "0000000000000000" & 
                           writeData(3 DOWNTO 2);    
                           writeData0_xhdl219 := "0000000000000000" & 
                           writeData(1 DOWNTO 0);    
                           CASE writeAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       wen_a71_xhdl146 := wen;    
                                       wen_a70_xhdl145 := wen;    
                                       wen_a69_xhdl144 := wen;    
                                       wen_a68_xhdl143 := wen;    
                                       wen_a67_xhdl142 := wen;    
                                       wen_a66_xhdl141 := wen;    
                                       wen_a65_xhdl140 := wen;    
                                       wen_a64_xhdl139 := wen;    
                                       wen_a63_xhdl138 := wen;    
                                       wen_a62_xhdl137 := wen;    
                                       wen_a61_xhdl136 := wen;    
                                       wen_a60_xhdl135 := wen;    
                                       wen_a59_xhdl134 := wen;    
                                       wen_a58_xhdl133 := wen;    
                                       wen_a57_xhdl132 := wen;    
                                       wen_a56_xhdl131 := wen;    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       wen_a71_xhdl146 := '0';    
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := wen;    
                                       wen_a54_xhdl129 := wen;    
                                       wen_a53_xhdl128 := wen;    
                                       wen_a52_xhdl127 := wen;    
                                       wen_a51_xhdl126 := wen;    
                                       wen_a50_xhdl125 := wen;    
                                       wen_a49_xhdl124 := wen;    
                                       wen_a48_xhdl123 := wen;    
                                       wen_a47_xhdl122 := wen;    
                                       wen_a46_xhdl121 := wen;    
                                       wen_a45_xhdl120 := wen;    
                                       wen_a44_xhdl119 := wen;    
                                       wen_a43_xhdl118 := wen;    
                                       wen_a42_xhdl117 := wen;    
                                       wen_a41_xhdl116 := wen;    
                                       wen_a40_xhdl115 := wen;    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       wen_a71_xhdl146 := '0';    
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := wen;    
                                       wen_a38_xhdl113 := wen;    
                                       wen_a37_xhdl112 := wen;    
                                       wen_a36_xhdl111 := wen;    
                                       wen_a35_xhdl110 := wen;    
                                       wen_a34_xhdl109 := wen;    
                                       wen_a33_xhdl108 := wen;    
                                       wen_a32_xhdl107 := wen;    
                                       wen_a31_xhdl106 := wen;    
                                       wen_a30_xhdl105 := wen;    
                                       wen_a29_xhdl104 := wen;    
                                       wen_a28_xhdl103 := wen;    
                                       wen_a27_xhdl102 := wen;    
                                       wen_a26_xhdl101 := wen;    
                                       wen_a25_xhdl100 := wen;    
                                       wen_a24_xhdl99 := wen;    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       wen_a71_xhdl146 := '0';    
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := wen;    
                                       wen_a22_xhdl97 := wen;    
                                       wen_a21_xhdl96 := wen;    
                                       wen_a20_xhdl95 := wen;    
                                       wen_a19_xhdl94 := wen;    
                                       wen_a18_xhdl93 := wen;    
                                       wen_a17_xhdl92 := wen;    
                                       wen_a16_xhdl91 := wen;    
                                       wen_a15_xhdl90 := wen;    
                                       wen_a14_xhdl89 := wen;    
                                       wen_a13_xhdl88 := wen;    
                                       wen_a12_xhdl87 := wen;    
                                       wen_a11_xhdl86 := wen;    
                                       wen_a10_xhdl85 := wen;    
                                       wen_a9_xhdl84 := wen;    
                                       wen_a8_xhdl83 := wen;    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" |
                                   "1000100" |
                                   "1000101" |
                                   "1000110" |
                                   "1000111" =>
                                       wen_a71_xhdl146 := '0';    
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := wen;    
                                       wen_a6_xhdl81 := wen;    
                                       wen_a5_xhdl80 := wen;    
                                       wen_a4_xhdl79 := wen;    
                                       wen_a3_xhdl78 := wen;    
                                       wen_a2_xhdl77 := wen;    
                                       wen_a1_xhdl76 := wen;    
                                       wen_a0_xhdl75 := wen;    
                              WHEN OTHERS  =>
                                       wen_a71_xhdl146 := '0';    
                                       wen_a70_xhdl145 := '0';    
                                       wen_a69_xhdl144 := '0';    
                                       wen_a68_xhdl143 := '0';    
                                       wen_a67_xhdl142 := '0';    
                                       wen_a66_xhdl141 := '0';    
                                       wen_a65_xhdl140 := '0';    
                                       wen_a64_xhdl139 := '0';    
                                       wen_a63_xhdl138 := '0';    
                                       wen_a62_xhdl137 := '0';    
                                       wen_a61_xhdl136 := '0';    
                                       wen_a60_xhdl135 := '0';    
                                       wen_a59_xhdl134 := '0';    
                                       wen_a58_xhdl133 := '0';    
                                       wen_a57_xhdl132 := '0';    
                                       wen_a56_xhdl131 := '0';    
                                       wen_a55_xhdl130 := '0';    
                                       wen_a54_xhdl129 := '0';    
                                       wen_a53_xhdl128 := '0';    
                                       wen_a52_xhdl127 := '0';    
                                       wen_a51_xhdl126 := '0';    
                                       wen_a50_xhdl125 := '0';    
                                       wen_a49_xhdl124 := '0';    
                                       wen_a48_xhdl123 := '0';    
                                       wen_a47_xhdl122 := '0';    
                                       wen_a46_xhdl121 := '0';    
                                       wen_a45_xhdl120 := '0';    
                                       wen_a44_xhdl119 := '0';    
                                       wen_a43_xhdl118 := '0';    
                                       wen_a42_xhdl117 := '0';    
                                       wen_a41_xhdl116 := '0';    
                                       wen_a40_xhdl115 := '0';    
                                       wen_a39_xhdl114 := '0';    
                                       wen_a38_xhdl113 := '0';    
                                       wen_a37_xhdl112 := '0';    
                                       wen_a36_xhdl111 := '0';    
                                       wen_a35_xhdl110 := '0';    
                                       wen_a34_xhdl109 := '0';    
                                       wen_a33_xhdl108 := '0';    
                                       wen_a32_xhdl107 := '0';    
                                       wen_a31_xhdl106 := '0';    
                                       wen_a30_xhdl105 := '0';    
                                       wen_a29_xhdl104 := '0';    
                                       wen_a28_xhdl103 := '0';    
                                       wen_a27_xhdl102 := '0';    
                                       wen_a26_xhdl101 := '0';    
                                       wen_a25_xhdl100 := '0';    
                                       wen_a24_xhdl99 := '0';    
                                       wen_a23_xhdl98 := '0';    
                                       wen_a22_xhdl97 := '0';    
                                       wen_a21_xhdl96 := '0';    
                                       wen_a20_xhdl95 := '0';    
                                       wen_a19_xhdl94 := '0';    
                                       wen_a18_xhdl93 := '0';    
                                       wen_a17_xhdl92 := '0';    
                                       wen_a16_xhdl91 := '0';    
                                       wen_a15_xhdl90 := '0';    
                                       wen_a14_xhdl89 := '0';    
                                       wen_a13_xhdl88 := '0';    
                                       wen_a12_xhdl87 := '0';    
                                       wen_a11_xhdl86 := '0';    
                                       wen_a10_xhdl85 := '0';    
                                       wen_a9_xhdl84 := '0';    
                                       wen_a8_xhdl83 := '0';    
                                       wen_a7_xhdl82 := '0';    
                                       wen_a6_xhdl81 := '0';    
                                       wen_a5_xhdl80 := '0';    
                                       wen_a4_xhdl79 := '0';    
                                       wen_a3_xhdl78 := '0';    
                                       wen_a2_xhdl77 := '0';    
                                       wen_a1_xhdl76 := '0';    
                                       wen_a0_xhdl75 := '0';    
                              
                              -- case: default
                              
                           END CASE;
                           -- case (writeAddr[11:6])
                           
                           CASE ckRdAddr(12 DOWNTO 6) IS
                              WHEN "0000000" |
                                   "0000001" |
                                   "0000010" |
                                   "0000011" |
                                   "0000100" |
                                   "0000101" |
                                   "0000110" |
                                   "0000111" |
                                   "0001000" |
                                   "0001001" |
                                   "0001010" |
                                   "0001011" |
                                   "0001100" |
                                   "0001101" |
                                   "0001110" |
                                   "0001111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData71(0)
                                       & readData70(0) & readData69(0) & 
                                       readData68(0) & readData67(0) & 
                                       readData66(0) & readData65(0) & 
                                       readData64(0) & readData63(0) & 
                                       readData62(0) & readData61(0) & 
                                       readData60(0) & readData59(0) & 
                                       readData58(0) & readData57(0) & 
                                       readData56(0);    
                              -- case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011, 7'b0000100, 7'b0000101,7'b0000110, 7'b0000111, 7'b0001000, 7'b0001001,...
                              
                              WHEN "0010000" |
                                   "0010001" |
                                   "0010010" |
                                   "0010011" |
                                   "0010100" |
                                   "0010101" |
                                   "0010110" |
                                   "0010111" |
                                   "0011000" |
                                   "0011001" |
                                   "0011010" |
                                   "0011011" |
                                   "0011100" |
                                   "0011101" |
                                   "0011110" |
                                   "0011111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData55(0)
                                       & readData54(0) & readData53(0) & 
                                       readData52(0) & readData51(0) & 
                                       readData50(0) & readData49(0) & 
                                       readData48(0) & readData47(0) & 
                                       readData46(0) & readData45(0) & 
                                       readData44(0) & readData43(0) & 
                                       readData42(0) & readData41(0) & 
                                       readData40(0);    
                              WHEN "0100000" |
                                   "0100001" |
                                   "0100010" |
                                   "0100011" |
                                   "0100100" |
                                   "0100101" |
                                   "0100110" |
                                   "0100111" |
                                   "0101000" |
                                   "0101001" |
                                   "0101010" |
                                   "0101011" |
                                   "0101100" |
                                   "0101101" |
                                   "0101110" |
                                   "0101111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData39(0)
                                       & readData38(0) & readData37(0) & 
                                       readData36(0) & readData35(0) & 
                                       readData34(0) & readData33(0) & 
                                       readData32(0) & readData31(0) & 
                                       readData30(0) & readData29(0) & 
                                       readData28(0) & readData27(0) & 
                                       readData26(0) & readData25(0) & 
                                       readData24(0);    
                              WHEN "0110000" |
                                   "0110001" |
                                   "0110010" |
                                   "0110011" |
                                   "0110100" |
                                   "0110101" |
                                   "0110110" |
                                   "0110111" |
                                   "0111000" |
                                   "0111001" |
                                   "0111010" |
                                   "0111011" |
                                   "0111100" |
                                   "0111101" |
                                   "0111110" |
                                   "0111111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData23(0)
                                       & readData22(0) & readData21(0) & 
                                       readData20(0) & readData19(0) & 
                                       readData18(0) & readData17(0) & 
                                       readData16(0) & readData15(0) & 
                                       readData14(0) & readData13(0) & 
                                       readData12(0) & readData11(0) & 
                                       readData10(0) & readData9(0) & 
                                       readData8(0);    
                              WHEN "1000000" |
                                   "1000001" |
                                   "1000010" |
                                   "1000011" |
                                   "1000100" |
                                   "1000101" |
                                   "1000110" |
                                   "1000111" =>
                                       readData_xhdl1_xhdl437_w16 := 
                                        readData7(1 
                                       DOWNTO 0) & readData6(1 DOWNTO 0) 
                                       & readData5(1 DOWNTO 0) & 
                                       readData4(1 DOWNTO 0) & 
                                       readData3(1 DOWNTO 0) & 
                                       readData2(1 DOWNTO 0) & 
                                       readData1(1 DOWNTO 0) & 
                                       readData0(1 DOWNTO 0);    
                              WHEN OTHERS  =>
                                       readData_xhdl1_xhdl437_w16 := (OTHERS 
                                       => '0');    
                              
                           END CASE;
                  WHEN OTHERS =>
                           NULL;
                  
               END CASE;
               -- case (USRAM_NUM_LOCATIONS_DWIDTH16)

      END IF;
      
      width0 <= width0_xhdl3;
      width1 <= width1_xhdl4;
      width2 <= width2_xhdl5;
      width3 <= width3_xhdl6;
      width4 <= width4_xhdl7;
      width5 <= width5_xhdl8;
      width6 <= width6_xhdl9;
      width7 <= width7_xhdl10;
      width8 <= width8_xhdl11;
      width9 <= width9_xhdl12;
      width10 <= width10_xhdl13;
      width11 <= width11_xhdl14;
      width12 <= width12_xhdl15;
      width13 <= width13_xhdl16;
      width14 <= width14_xhdl17;
      width15 <= width15_xhdl18;
      width16 <= width16_xhdl19;
      width17 <= width17_xhdl20;
      width18 <= width18_xhdl21;
      width19 <= width19_xhdl22;
      width20 <= width20_xhdl23;
      width21 <= width21_xhdl24;
      width22 <= width22_xhdl25;
      width23 <= width23_xhdl26;
      width24 <= width24_xhdl27;
      width25 <= width25_xhdl28;
      width26 <= width26_xhdl29;
      width27 <= width27_xhdl30;
      width28 <= width28_xhdl31;
      width29 <= width29_xhdl32;
      width30 <= width30_xhdl33;
      width31 <= width31_xhdl34;
      width32 <= width32_xhdl35;
      width33 <= width33_xhdl36;
      width34 <= width34_xhdl37;
      width35 <= width35_xhdl38;
      width36 <= width36_xhdl39;
      width37 <= width37_xhdl40;
      width38 <= width38_xhdl41;
      width39 <= width39_xhdl42;
      width40 <= width40_xhdl43;
      width41 <= width41_xhdl44;
      width42 <= width42_xhdl45;
      width43 <= width43_xhdl46;
      width44 <= width44_xhdl47;
      width45 <= width45_xhdl48;
      width46 <= width46_xhdl49;
      width47 <= width47_xhdl50;
      width48 <= width48_xhdl51;
      width49 <= width49_xhdl52;
      width50 <= width50_xhdl53;
      width51 <= width51_xhdl54;
      width52 <= width52_xhdl55;
      width53 <= width53_xhdl56;
      width54 <= width54_xhdl57;
      width55 <= width55_xhdl58;
      width56 <= width56_xhdl59;
      width57 <= width57_xhdl60;
      width58 <= width58_xhdl61;
      width59 <= width59_xhdl62;
      width60 <= width60_xhdl63;
      width61 <= width61_xhdl64;
      width62 <= width62_xhdl65;
      width63 <= width63_xhdl66;
      width64 <= width64_xhdl67;
      width65 <= width65_xhdl68;
      width66 <= width66_xhdl69;
      width67 <= width67_xhdl70;
      width68 <= width68_xhdl71;
      width69 <= width69_xhdl72;
      width70 <= width70_xhdl73;
      width71 <= width71_xhdl74;
      wen_a0 <= wen_a0_xhdl75;
      wen_a1 <= wen_a1_xhdl76;
      wen_a2 <= wen_a2_xhdl77;
      wen_a3 <= wen_a3_xhdl78;
      wen_a4 <= wen_a4_xhdl79;
      wen_a5 <= wen_a5_xhdl80;
      wen_a6 <= wen_a6_xhdl81;
      wen_a7 <= wen_a7_xhdl82;
      wen_a8 <= wen_a8_xhdl83;
      wen_a9 <= wen_a9_xhdl84;
      wen_a10 <= wen_a10_xhdl85;
      wen_a11 <= wen_a11_xhdl86;
      wen_a12 <= wen_a12_xhdl87;
      wen_a13 <= wen_a13_xhdl88;
      wen_a14 <= wen_a14_xhdl89;
      wen_a15 <= wen_a15_xhdl90;
      wen_a16 <= wen_a16_xhdl91;
      wen_a17 <= wen_a17_xhdl92;
      wen_a18 <= wen_a18_xhdl93;
      wen_a19 <= wen_a19_xhdl94;
      wen_a20 <= wen_a20_xhdl95;
      wen_a21 <= wen_a21_xhdl96;
      wen_a22 <= wen_a22_xhdl97;
      wen_a23 <= wen_a23_xhdl98;
      wen_a24 <= wen_a24_xhdl99;
      wen_a25 <= wen_a25_xhdl100;
      wen_a26 <= wen_a26_xhdl101;
      wen_a27 <= wen_a27_xhdl102;
      wen_a28 <= wen_a28_xhdl103;
      wen_a29 <= wen_a29_xhdl104;
      wen_a30 <= wen_a30_xhdl105;
      wen_a31 <= wen_a31_xhdl106;
      wen_a32 <= wen_a32_xhdl107;
      wen_a33 <= wen_a33_xhdl108;
      wen_a34 <= wen_a34_xhdl109;
      wen_a35 <= wen_a35_xhdl110;
      wen_a36 <= wen_a36_xhdl111;
      wen_a37 <= wen_a37_xhdl112;
      wen_a38 <= wen_a38_xhdl113;
      wen_a39 <= wen_a39_xhdl114;
      wen_a40 <= wen_a40_xhdl115;
      wen_a41 <= wen_a41_xhdl116;
      wen_a42 <= wen_a42_xhdl117;
      wen_a43 <= wen_a43_xhdl118;
      wen_a44 <= wen_a44_xhdl119;
      wen_a45 <= wen_a45_xhdl120;
      wen_a46 <= wen_a46_xhdl121;
      wen_a47 <= wen_a47_xhdl122;
      wen_a48 <= wen_a48_xhdl123;
      wen_a49 <= wen_a49_xhdl124;
      wen_a50 <= wen_a50_xhdl125;
      wen_a51 <= wen_a51_xhdl126;
      wen_a52 <= wen_a52_xhdl127;
      wen_a53 <= wen_a53_xhdl128;
      wen_a54 <= wen_a54_xhdl129;
      wen_a55 <= wen_a55_xhdl130;
      wen_a56 <= wen_a56_xhdl131;
      wen_a57 <= wen_a57_xhdl132;
      wen_a58 <= wen_a58_xhdl133;
      wen_a59 <= wen_a59_xhdl134;
      wen_a60 <= wen_a60_xhdl135;
      wen_a61 <= wen_a61_xhdl136;
      wen_a62 <= wen_a62_xhdl137;
      wen_a63 <= wen_a63_xhdl138;
      wen_a64 <= wen_a64_xhdl139;
      wen_a65 <= wen_a65_xhdl140;
      wen_a66 <= wen_a66_xhdl141;
      wen_a67 <= wen_a67_xhdl142;
      wen_a68 <= wen_a68_xhdl143;
      wen_a69 <= wen_a69_xhdl144;
      wen_a70 <= wen_a70_xhdl145;
      wen_a71 <= wen_a71_xhdl146;
      wen_b0 <= wen_b0_xhdl147;
      wen_b1 <= wen_b1_xhdl148;
      wen_b2 <= wen_b2_xhdl149;
      wen_b3 <= wen_b3_xhdl150;
      wen_b4 <= wen_b4_xhdl151;
      wen_b5 <= wen_b5_xhdl152;
      wen_b6 <= wen_b6_xhdl153;
      wen_b7 <= wen_b7_xhdl154;
      wen_b8 <= wen_b8_xhdl155;
      wen_b9 <= wen_b9_xhdl156;
      wen_b10 <= wen_b10_xhdl157;
      wen_b11 <= wen_b11_xhdl158;
      wen_b12 <= wen_b12_xhdl159;
      wen_b13 <= wen_b13_xhdl160;
      wen_b14 <= wen_b14_xhdl161;
      wen_b15 <= wen_b15_xhdl162;
      wen_b16 <= wen_b16_xhdl163;
      wen_b17 <= wen_b17_xhdl164;
      wen_b18 <= wen_b18_xhdl165;
      wen_b19 <= wen_b19_xhdl166;
      wen_b20 <= wen_b20_xhdl167;
      wen_b21 <= wen_b21_xhdl168;
      wen_b22 <= wen_b22_xhdl169;
      wen_b23 <= wen_b23_xhdl170;
      wen_b24 <= wen_b24_xhdl171;
      wen_b25 <= wen_b25_xhdl172;
      wen_b26 <= wen_b26_xhdl173;
      wen_b27 <= wen_b27_xhdl174;
      wen_b28 <= wen_b28_xhdl175;
      wen_b29 <= wen_b29_xhdl176;
      wen_b30 <= wen_b30_xhdl177;
      wen_b31 <= wen_b31_xhdl178;
      wen_b32 <= wen_b32_xhdl179;
      wen_b33 <= wen_b33_xhdl180;
      wen_b34 <= wen_b34_xhdl181;
      wen_b35 <= wen_b35_xhdl182;
      wen_b36 <= wen_b36_xhdl183;
      wen_b37 <= wen_b37_xhdl184;
      wen_b38 <= wen_b38_xhdl185;
      wen_b39 <= wen_b39_xhdl186;
      wen_b40 <= wen_b40_xhdl187;
      wen_b41 <= wen_b41_xhdl188;
      wen_b42 <= wen_b42_xhdl189;
      wen_b43 <= wen_b43_xhdl190;
      wen_b44 <= wen_b44_xhdl191;
      wen_b45 <= wen_b45_xhdl192;
      wen_b46 <= wen_b46_xhdl193;
      wen_b47 <= wen_b47_xhdl194;
      wen_b48 <= wen_b48_xhdl195;
      wen_b49 <= wen_b49_xhdl196;
      wen_b50 <= wen_b50_xhdl197;
      wen_b51 <= wen_b51_xhdl198;
      wen_b52 <= wen_b52_xhdl199;
      wen_b53 <= wen_b53_xhdl200;
      wen_b54 <= wen_b54_xhdl201;
      wen_b55 <= wen_b55_xhdl202;
      wen_b56 <= wen_b56_xhdl203;
      wen_b57 <= wen_b57_xhdl204;
      wen_b58 <= wen_b58_xhdl205;
      wen_b59 <= wen_b59_xhdl206;
      wen_b60 <= wen_b60_xhdl207;
      wen_b61 <= wen_b61_xhdl208;
      wen_b62 <= wen_b62_xhdl209;
      wen_b63 <= wen_b63_xhdl210;
      wen_b64 <= wen_b64_xhdl211;
      wen_b65 <= wen_b65_xhdl212;
      wen_b66 <= wen_b66_xhdl213;
      wen_b67 <= wen_b67_xhdl214;
      wen_b68 <= wen_b68_xhdl215;
      wen_b69 <= wen_b69_xhdl216;
      wen_b70 <= wen_b70_xhdl217;
      wen_b71 <= wen_b71_xhdl218;
      writeData0 <= writeData0_xhdl219;
      writeData1 <= writeData1_xhdl220;
      writeData2 <= writeData2_xhdl221;
      writeData3 <= writeData3_xhdl222;
      writeData4 <= writeData4_xhdl223;
      writeData5 <= writeData5_xhdl224;
      writeData6 <= writeData6_xhdl225;
      writeData7 <= writeData7_xhdl226;
      writeData8 <= writeData8_xhdl227;
      writeData9 <= writeData9_xhdl228;
      writeData10 <= writeData10_xhdl229;
      writeData11 <= writeData11_xhdl230;
      writeData12 <= writeData12_xhdl231;
      writeData13 <= writeData13_xhdl232;
      writeData14 <= writeData14_xhdl233;
      writeData15 <= writeData15_xhdl234;
      writeData16 <= writeData16_xhdl235;
      writeData17 <= writeData17_xhdl236;
      writeData18 <= writeData18_xhdl237;
      writeData19 <= writeData19_xhdl238;
      writeData20 <= writeData20_xhdl239;
      writeData21 <= writeData21_xhdl240;
      writeData22 <= writeData22_xhdl241;
      writeData23 <= writeData23_xhdl242;
      writeData24 <= writeData24_xhdl243;
      writeData25 <= writeData25_xhdl244;
      writeData26 <= writeData26_xhdl245;
      writeData27 <= writeData27_xhdl246;
      writeData28 <= writeData28_xhdl247;
      writeData29 <= writeData29_xhdl248;
      writeData30 <= writeData30_xhdl249;
      writeData31 <= writeData31_xhdl250;
      writeData32 <= writeData32_xhdl251;
      writeData33 <= writeData33_xhdl252;
      writeData34 <= writeData34_xhdl253;
      writeData35 <= writeData35_xhdl254;
      writeData36 <= writeData36_xhdl255;
      writeData37 <= writeData37_xhdl256;
      writeData38 <= writeData38_xhdl257;
      writeData39 <= writeData39_xhdl258;
      writeData40 <= writeData40_xhdl259;
      writeData41 <= writeData41_xhdl260;
      writeData42 <= writeData42_xhdl261;
      writeData43 <= writeData43_xhdl262;
      writeData44 <= writeData44_xhdl263;
      writeData45 <= writeData45_xhdl264;
      writeData46 <= writeData46_xhdl265;
      writeData47 <= writeData47_xhdl266;
      writeData48 <= writeData48_xhdl267;
      writeData49 <= writeData49_xhdl268;
      writeData50 <= writeData50_xhdl269;
      writeData51 <= writeData51_xhdl270;
      writeData52 <= writeData52_xhdl271;
      writeData53 <= writeData53_xhdl272;
      writeData54 <= writeData54_xhdl273;
      writeData55 <= writeData55_xhdl274;
      writeData56 <= writeData56_xhdl275;
      writeData57 <= writeData57_xhdl276;
      writeData58 <= writeData58_xhdl277;
      writeData59 <= writeData59_xhdl278;
      writeData60 <= writeData60_xhdl279;
      writeData61 <= writeData61_xhdl280;
      writeData62 <= writeData62_xhdl281;
      writeData63 <= writeData63_xhdl282;
      writeData64 <= writeData64_xhdl283;
      writeData65 <= writeData65_xhdl284;
      writeData66 <= writeData66_xhdl285;
      writeData67 <= writeData67_xhdl286;
      writeData68 <= writeData68_xhdl287;
      writeData69 <= writeData69_xhdl288;
      writeData70 <= writeData70_xhdl289;
      writeData71 <= writeData71_xhdl290;
      writeAddr0 <= writeAddr0_xhdl291;
      writeAddr1 <= writeAddr1_xhdl292;
      writeAddr2 <= writeAddr2_xhdl293;
      writeAddr3 <= writeAddr3_xhdl294;
      writeAddr4 <= writeAddr4_xhdl295;
      writeAddr5 <= writeAddr5_xhdl296;
      writeAddr6 <= writeAddr6_xhdl297;
      writeAddr7 <= writeAddr7_xhdl298;
      writeAddr8 <= writeAddr8_xhdl299;
      writeAddr9 <= writeAddr9_xhdl300;
      writeAddr10 <= writeAddr10_xhdl301;
      writeAddr11 <= writeAddr11_xhdl302;
      writeAddr12 <= writeAddr12_xhdl303;
      writeAddr13 <= writeAddr13_xhdl304;
      writeAddr14 <= writeAddr14_xhdl305;
      writeAddr15 <= writeAddr15_xhdl306;
      writeAddr16 <= writeAddr16_xhdl307;
      writeAddr17 <= writeAddr17_xhdl308;
      writeAddr18 <= writeAddr18_xhdl309;
      writeAddr19 <= writeAddr19_xhdl310;
      writeAddr20 <= writeAddr20_xhdl311;
      writeAddr21 <= writeAddr21_xhdl312;
      writeAddr22 <= writeAddr22_xhdl313;
      writeAddr23 <= writeAddr23_xhdl314;
      writeAddr24 <= writeAddr24_xhdl315;
      writeAddr25 <= writeAddr25_xhdl316;
      writeAddr26 <= writeAddr26_xhdl317;
      writeAddr27 <= writeAddr27_xhdl318;
      writeAddr28 <= writeAddr28_xhdl319;
      writeAddr29 <= writeAddr29_xhdl320;
      writeAddr30 <= writeAddr30_xhdl321;
      writeAddr31 <= writeAddr31_xhdl322;
      writeAddr32 <= writeAddr32_xhdl323;
      writeAddr33 <= writeAddr33_xhdl324;
      writeAddr34 <= writeAddr34_xhdl325;
      writeAddr35 <= writeAddr35_xhdl326;
      writeAddr36 <= writeAddr36_xhdl327;
      writeAddr37 <= writeAddr37_xhdl328;
      writeAddr38 <= writeAddr38_xhdl329;
      writeAddr39 <= writeAddr39_xhdl330;
      writeAddr40 <= writeAddr40_xhdl331;
      writeAddr41 <= writeAddr41_xhdl332;
      writeAddr42 <= writeAddr42_xhdl333;
      writeAddr43 <= writeAddr43_xhdl334;
      writeAddr44 <= writeAddr44_xhdl335;
      writeAddr45 <= writeAddr45_xhdl336;
      writeAddr46 <= writeAddr46_xhdl337;
      writeAddr47 <= writeAddr47_xhdl338;
      writeAddr48 <= writeAddr48_xhdl339;
      writeAddr49 <= writeAddr49_xhdl340;
      writeAddr50 <= writeAddr50_xhdl341;
      writeAddr51 <= writeAddr51_xhdl342;
      writeAddr52 <= writeAddr52_xhdl343;
      writeAddr53 <= writeAddr53_xhdl344;
      writeAddr54 <= writeAddr54_xhdl345;
      writeAddr55 <= writeAddr55_xhdl346;
      writeAddr56 <= writeAddr56_xhdl347;
      writeAddr57 <= writeAddr57_xhdl348;
      writeAddr58 <= writeAddr58_xhdl349;
      writeAddr59 <= writeAddr59_xhdl350;
      writeAddr60 <= writeAddr60_xhdl351;
      writeAddr61 <= writeAddr61_xhdl352;
      writeAddr62 <= writeAddr62_xhdl353;
      writeAddr63 <= writeAddr63_xhdl354;
      writeAddr64 <= writeAddr64_xhdl355;
      writeAddr65 <= writeAddr65_xhdl356;
      writeAddr66 <= writeAddr66_xhdl357;
      writeAddr67 <= writeAddr67_xhdl358;
      writeAddr68 <= writeAddr68_xhdl359;
      writeAddr69 <= writeAddr69_xhdl360;
      writeAddr70 <= writeAddr70_xhdl361;
      writeAddr71 <= writeAddr71_xhdl362;
      readAddr0 <= readAddr0_xhdl363;
      readAddr1 <= readAddr1_xhdl364;
      readAddr2 <= readAddr2_xhdl365;
      readAddr3 <= readAddr3_xhdl366;
      readAddr4 <= readAddr4_xhdl367;
      readAddr5 <= readAddr5_xhdl368;
      readAddr6 <= readAddr6_xhdl369;
      readAddr7 <= readAddr7_xhdl370;
      readAddr8 <= readAddr8_xhdl371;
      readAddr9 <= readAddr9_xhdl372;
      readAddr10 <= readAddr10_xhdl373;
      readAddr11 <= readAddr11_xhdl374;
      readAddr12 <= readAddr12_xhdl375;
      readAddr13 <= readAddr13_xhdl376;
      readAddr14 <= readAddr14_xhdl377;
      readAddr15 <= readAddr15_xhdl378;
      readAddr16 <= readAddr16_xhdl379;
      readAddr17 <= readAddr17_xhdl380;
      readAddr18 <= readAddr18_xhdl381;
      readAddr19 <= readAddr19_xhdl382;
      readAddr20 <= readAddr20_xhdl383;
      readAddr21 <= readAddr21_xhdl384;
      readAddr22 <= readAddr22_xhdl385;
      readAddr23 <= readAddr23_xhdl386;
      readAddr24 <= readAddr24_xhdl387;
      readAddr25 <= readAddr25_xhdl388;
      readAddr26 <= readAddr26_xhdl389;
      readAddr27 <= readAddr27_xhdl390;
      readAddr28 <= readAddr28_xhdl391;
      readAddr29 <= readAddr29_xhdl392;
      readAddr30 <= readAddr30_xhdl393;
      readAddr31 <= readAddr31_xhdl394;
      readAddr32 <= readAddr32_xhdl395;
      readAddr33 <= readAddr33_xhdl396;
      readAddr34 <= readAddr34_xhdl397;
      readAddr35 <= readAddr35_xhdl398;
      readAddr36 <= readAddr36_xhdl399;
      readAddr37 <= readAddr37_xhdl400;
      readAddr38 <= readAddr38_xhdl401;
      readAddr39 <= readAddr39_xhdl402;
      readAddr40 <= readAddr40_xhdl403;
      readAddr41 <= readAddr41_xhdl404;
      readAddr42 <= readAddr42_xhdl405;
      readAddr43 <= readAddr43_xhdl406;
      readAddr44 <= readAddr44_xhdl407;
      readAddr45 <= readAddr45_xhdl408;
      readAddr46 <= readAddr46_xhdl409;
      readAddr47 <= readAddr47_xhdl410;
      readAddr48 <= readAddr48_xhdl411;
      readAddr49 <= readAddr49_xhdl412;
      readAddr50 <= readAddr50_xhdl413;
      readAddr51 <= readAddr51_xhdl414;
      readAddr52 <= readAddr52_xhdl415;
      readAddr53 <= readAddr53_xhdl416;
      readAddr54 <= readAddr54_xhdl417;
      readAddr55 <= readAddr55_xhdl418;
      readAddr56 <= readAddr56_xhdl419;
      readAddr57 <= readAddr57_xhdl420;
      readAddr58 <= readAddr58_xhdl421;
      readAddr59 <= readAddr59_xhdl422;
      readAddr60 <= readAddr60_xhdl423;
      readAddr61 <= readAddr61_xhdl424;
      readAddr62 <= readAddr62_xhdl425;
      readAddr63 <= readAddr63_xhdl426;
      readAddr64 <= readAddr64_xhdl427;
      readAddr65 <= readAddr65_xhdl428;
      readAddr66 <= readAddr66_xhdl429;
      readAddr67 <= readAddr67_xhdl430;
      readAddr68 <= readAddr68_xhdl431;
      readAddr69 <= readAddr69_xhdl432;
      readAddr70 <= readAddr70_xhdl433;
      readAddr71 <= readAddr71_xhdl434;
      ablk <= ablk_xhdl435 after 1ns;
      bblk <= bblk_xhdl436 after 1ns;
      cblk <= cblk_xhdl437;

      readData_xhdl1 <= readData_xhdl1_xhdl437_w16;

   END PROCESS;
   
   -- always @ (*)
   ------------------------------------------------------------------------------------------
   -- RAM64x18 blocks
   ------------------------------------------------------------------------------------------
   block_71 : RAM64x18 
      PORT MAP (
         A_DOUT => readData71,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr71,
         B_ADDR => readAddr71,
         A_WIDTH => width71,
         B_WIDTH => width71,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr71,
         C_DIN => writeData71,
         C_WEN => wen_a71,
         C_BLK => cblk,
         C_WIDTH => width71,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_71);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_70 : RAM64x18 
      PORT MAP (
         A_DOUT => readData70,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr70,
         B_ADDR => readAddr70,
         A_WIDTH => width70,
         B_WIDTH => width70,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr70,
         C_DIN => writeData70,
         C_WEN => wen_a70,
         C_BLK => cblk,
         C_WIDTH => width70,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_70);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_69 : RAM64x18 
      PORT MAP (
         A_DOUT => readData69,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr69,
         B_ADDR => readAddr69,
         A_WIDTH => width69,
         B_WIDTH => width69,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr69,
         C_DIN => writeData69,
         C_WEN => wen_a69,
         C_BLK => cblk,
         C_WIDTH => width69,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_69);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_68 : RAM64x18 
      PORT MAP (
         A_DOUT => readData68,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr68,
         B_ADDR => readAddr68,
         A_WIDTH => width68,
         B_WIDTH => width68,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr68,
         C_DIN => writeData68,
         C_WEN => wen_a68,
         C_BLK => cblk,
         C_WIDTH => width68,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_68);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_67 : RAM64x18 
      PORT MAP (
         A_DOUT => readData67,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr67,
         B_ADDR => readAddr67,
         A_WIDTH => width67,
         B_WIDTH => width67,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr67,
         C_DIN => writeData67,
         C_WEN => wen_a67,
         C_BLK => cblk,
         C_WIDTH => width67,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_67);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_66 : RAM64x18 
      PORT MAP (
         A_DOUT => readData66,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr66,
         B_ADDR => readAddr66,
         A_WIDTH => width66,
         B_WIDTH => width66,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr66,
         C_DIN => writeData66,
         C_WEN => wen_a66,
         C_BLK => cblk,
         C_WIDTH => width66,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_66);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_65 : RAM64x18 
      PORT MAP (
         A_DOUT => readData65,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr65,
         B_ADDR => readAddr65,
         A_WIDTH => width65,
         B_WIDTH => width65,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr65,
         C_DIN => writeData65,
         C_WEN => wen_a65,
         C_BLK => cblk,
         C_WIDTH => width65,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_65);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_64 : RAM64x18 
      PORT MAP (
         A_DOUT => readData64,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr64,
         B_ADDR => readAddr64,
         A_WIDTH => width64,
         B_WIDTH => width64,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr64,
         C_DIN => writeData64,
         C_WEN => wen_a64,
         C_BLK => cblk,
         C_WIDTH => width64,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_64);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_63 : RAM64x18 
      PORT MAP (
         A_DOUT => readData63,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr63,
         B_ADDR => readAddr63,
         A_WIDTH => width63,
         B_WIDTH => width63,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr63,
         C_DIN => writeData63,
         C_WEN => wen_a63,
         C_BLK => cblk,
         C_WIDTH => width63,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_63);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_62 : RAM64x18 
      PORT MAP (
         A_DOUT => readData62,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr62,
         B_ADDR => readAddr62,
         A_WIDTH => width62,
         B_WIDTH => width62,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr62,
         C_DIN => writeData62,
         C_WEN => wen_a62,
         C_BLK => cblk,
         C_WIDTH => width62,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_62);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_61 : RAM64x18 
      PORT MAP (
         A_DOUT => readData61,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr61,
         B_ADDR => readAddr61,
         A_WIDTH => width61,
         B_WIDTH => width61,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr61,
         C_DIN => writeData61,
         C_WEN => wen_a61,
         C_BLK => cblk,
         C_WIDTH => width61,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_61);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_60 : RAM64x18 
      PORT MAP (
         A_DOUT => readData60,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr60,
         B_ADDR => readAddr60,
         A_WIDTH => width60,
         B_WIDTH => width60,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr60,
         C_DIN => writeData60,
         C_WEN => wen_a60,
         C_BLK => cblk,
         C_WIDTH => width60,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_60);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_59 : RAM64x18 
      PORT MAP (
         A_DOUT => readData59,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr59,
         B_ADDR => readAddr59,
         A_WIDTH => width59,
         B_WIDTH => width59,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr59,
         C_DIN => writeData59,
         C_WEN => wen_a59,
         C_BLK => cblk,
         C_WIDTH => width59,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_59);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_58 : RAM64x18 
      PORT MAP (
         A_DOUT => readData58,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr58,
         B_ADDR => readAddr58,
         A_WIDTH => width58,
         B_WIDTH => width58,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr58,
         C_DIN => writeData58,
         C_WEN => wen_a58,
         C_BLK => cblk,
         C_WIDTH => width58,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_58);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_57 : RAM64x18 
      PORT MAP (
         A_DOUT => readData57,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr57,
         B_ADDR => readAddr57,
         A_WIDTH => width57,
         B_WIDTH => width57,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr57,
         C_DIN => writeData57,
         C_WEN => wen_a57,
         C_BLK => cblk,
         C_WIDTH => width57,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_57);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_56 : RAM64x18 
      PORT MAP (
         A_DOUT => readData56,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr56,
         B_ADDR => readAddr56,
         A_WIDTH => width56,
         B_WIDTH => width56,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr56,
         C_DIN => writeData56,
         C_WEN => wen_a56,
         C_BLK => cblk,
         C_WIDTH => width56,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_56);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_55 : RAM64x18 
      PORT MAP (
         A_DOUT => readData55,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr55,
         B_ADDR => readAddr55,
         A_WIDTH => width55,
         B_WIDTH => width55,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr55,
         C_DIN => writeData55,
         C_WEN => wen_a55,
         C_BLK => cblk,
         C_WIDTH => width55,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_55);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_54 : RAM64x18 
      PORT MAP (
         A_DOUT => readData54,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr54,
         B_ADDR => readAddr54,
         A_WIDTH => width54,
         B_WIDTH => width54,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr54,
         C_DIN => writeData54,
         C_WEN => wen_a54,
         C_BLK => cblk,
         C_WIDTH => width54,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_54);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_53 : RAM64x18 
      PORT MAP (
         A_DOUT => readData53,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr53,
         B_ADDR => readAddr53,
         A_WIDTH => width53,
         B_WIDTH => width53,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr53,
         C_DIN => writeData53,
         C_WEN => wen_a53,
         C_BLK => cblk,
         C_WIDTH => width53,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_53);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_52 : RAM64x18 
      PORT MAP (
         A_DOUT => readData52,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr52,
         B_ADDR => readAddr52,
         A_WIDTH => width52,
         B_WIDTH => width52,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr52,
         C_DIN => writeData52,
         C_WEN => wen_a52,
         C_BLK => cblk,
         C_WIDTH => width52,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_52);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_51 : RAM64x18 
      PORT MAP (
         A_DOUT => readData51,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr51,
         B_ADDR => readAddr51,
         A_WIDTH => width51,
         B_WIDTH => width51,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr51,
         C_DIN => writeData51,
         C_WEN => wen_a51,
         C_BLK => cblk,
         C_WIDTH => width51,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_51);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_50 : RAM64x18 
      PORT MAP (
         A_DOUT => readData50,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr50,
         B_ADDR => readAddr50,
         A_WIDTH => width50,
         B_WIDTH => width50,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr50,
         C_DIN => writeData50,
         C_WEN => wen_a50,
         C_BLK => cblk,
         C_WIDTH => width50,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_50);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_49 : RAM64x18 
      PORT MAP (
         A_DOUT => readData49,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr49,
         B_ADDR => readAddr49,
         A_WIDTH => width49,
         B_WIDTH => width49,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr49,
         C_DIN => writeData49,
         C_WEN => wen_a49,
         C_BLK => cblk,
         C_WIDTH => width49,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_49);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_48 : RAM64x18 
      PORT MAP (
         A_DOUT => readData48,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr48,
         B_ADDR => readAddr48,
         A_WIDTH => width48,
         B_WIDTH => width48,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr48,
         C_DIN => writeData48,
         C_WEN => wen_a48,
         C_BLK => cblk,
         C_WIDTH => width48,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_48);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_47 : RAM64x18 
      PORT MAP (
         A_DOUT => readData47,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr47,
         B_ADDR => readAddr47,
         A_WIDTH => width47,
         B_WIDTH => width47,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr47,
         C_DIN => writeData47,
         C_WEN => wen_a47,
         C_BLK => cblk,
         C_WIDTH => width47,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_47);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_46 : RAM64x18 
      PORT MAP (
         A_DOUT => readData46,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr46,
         B_ADDR => readAddr46,
         A_WIDTH => width46,
         B_WIDTH => width46,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr46,
         C_DIN => writeData46,
         C_WEN => wen_a46,
         C_BLK => cblk,
         C_WIDTH => width46,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_46);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_45 : RAM64x18 
      PORT MAP (
         A_DOUT => readData45,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr45,
         B_ADDR => readAddr45,
         A_WIDTH => width45,
         B_WIDTH => width45,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr45,
         C_DIN => writeData45,
         C_WEN => wen_a45,
         C_BLK => cblk,
         C_WIDTH => width45,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_45);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_44 : RAM64x18 
      PORT MAP (
         A_DOUT => readData44,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr44,
         B_ADDR => readAddr44,
         A_WIDTH => width44,
         B_WIDTH => width44,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr44,
         C_DIN => writeData44,
         C_WEN => wen_a44,
         C_BLK => cblk,
         C_WIDTH => width44,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_44);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_43 : RAM64x18 
      PORT MAP (
         A_DOUT => readData43,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr43,
         B_ADDR => readAddr43,
         A_WIDTH => width43,
         B_WIDTH => width43,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr43,
         C_DIN => writeData43,
         C_WEN => wen_a43,
         C_BLK => cblk,
         C_WIDTH => width43,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_43);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_42 : RAM64x18 
      PORT MAP (
         A_DOUT => readData42,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr42,
         B_ADDR => readAddr42,
         A_WIDTH => width42,
         B_WIDTH => width42,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr42,
         C_DIN => writeData42,
         C_WEN => wen_a42,
         C_BLK => cblk,
         C_WIDTH => width42,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_42);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_41 : RAM64x18 
      PORT MAP (
         A_DOUT => readData41,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr41,
         B_ADDR => readAddr41,
         A_WIDTH => width41,
         B_WIDTH => width41,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr41,
         C_DIN => writeData41,
         C_WEN => wen_a41,
         C_BLK => cblk,
         C_WIDTH => width41,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_41);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_40 : RAM64x18 
      PORT MAP (
         A_DOUT => readData40,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr40,
         B_ADDR => readAddr40,
         A_WIDTH => width40,
         B_WIDTH => width40,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr40,
         C_DIN => writeData40,
         C_WEN => wen_a40,
         C_BLK => cblk,
         C_WIDTH => width40,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_40);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_39 : RAM64x18 
      PORT MAP (
         A_DOUT => readData39,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr39,
         B_ADDR => readAddr39,
         A_WIDTH => width39,
         B_WIDTH => width39,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr39,
         C_DIN => writeData39,
         C_WEN => wen_a39,
         C_BLK => cblk,
         C_WIDTH => width39,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_39);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_38 : RAM64x18 
      PORT MAP (
         A_DOUT => readData38,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr38,
         B_ADDR => readAddr38,
         A_WIDTH => width38,
         B_WIDTH => width38,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr38,
         C_DIN => writeData38,
         C_WEN => wen_a38,
         C_BLK => cblk,
         C_WIDTH => width38,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_38);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_37 : RAM64x18 
      PORT MAP (
         A_DOUT => readData37,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr37,
         B_ADDR => readAddr37,
         A_WIDTH => width37,
         B_WIDTH => width37,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr37,
         C_DIN => writeData37,
         C_WEN => wen_a37,
         C_BLK => cblk,
         C_WIDTH => width37,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_37);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_36 : RAM64x18 
      PORT MAP (
         A_DOUT => readData36,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr36,
         B_ADDR => readAddr36,
         A_WIDTH => width36,
         B_WIDTH => width36,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr36,
         C_DIN => writeData36,
         C_WEN => wen_a36,
         C_BLK => cblk,
         C_WIDTH => width36,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_36);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_35 : RAM64x18 
      PORT MAP (
         A_DOUT => readData35,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr35,
         B_ADDR => readAddr35,
         A_WIDTH => width35,
         B_WIDTH => width35,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr35,
         C_DIN => writeData35,
         C_WEN => wen_a35,
         C_BLK => cblk,
         C_WIDTH => width35,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_35);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_34 : RAM64x18 
      PORT MAP (
         A_DOUT => readData34,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr34,
         B_ADDR => readAddr34,
         A_WIDTH => width34,
         B_WIDTH => width34,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr34,
         C_DIN => writeData34,
         C_WEN => wen_a34,
         C_BLK => cblk,
         C_WIDTH => width34,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_34);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_33 : RAM64x18 
      PORT MAP (
         A_DOUT => readData33,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr33,
         B_ADDR => readAddr33,
         A_WIDTH => width33,
         B_WIDTH => width33,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr33,
         C_DIN => writeData33,
         C_WEN => wen_a33,
         C_BLK => cblk,
         C_WIDTH => width33,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_33);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_32 : RAM64x18 
      PORT MAP (
         A_DOUT => readData32,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr32,
         B_ADDR => readAddr32,
         A_WIDTH => width32,
         B_WIDTH => width32,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr32,
         C_DIN => writeData32,
         C_WEN => wen_a32,
         C_BLK => cblk,
         C_WIDTH => width32,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_32);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_31 : RAM64x18 
      PORT MAP (
         A_DOUT => readData31,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr31,
         B_ADDR => readAddr31,
         A_WIDTH => width31,
         B_WIDTH => width31,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr31,
         C_DIN => writeData31,
         C_WEN => wen_a31,
         C_BLK => cblk,
         C_WIDTH => width31,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_31);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_30 : RAM64x18 
      PORT MAP (
         A_DOUT => readData30,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr30,
         B_ADDR => readAddr30,
         A_WIDTH => width30,
         B_WIDTH => width30,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr30,
         C_DIN => writeData30,
         C_WEN => wen_a30,
         C_BLK => cblk,
         C_WIDTH => width30,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_30);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_29 : RAM64x18 
      PORT MAP (
         A_DOUT => readData29,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr29,
         B_ADDR => readAddr29,
         A_WIDTH => width29,
         B_WIDTH => width29,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr29,
         C_DIN => writeData29,
         C_WEN => wen_a29,
         C_BLK => cblk,
         C_WIDTH => width29,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_29);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_28 : RAM64x18 
      PORT MAP (
         A_DOUT => readData28,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr28,
         B_ADDR => readAddr28,
         A_WIDTH => width28,
         B_WIDTH => width28,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr28,
         C_DIN => writeData28,
         C_WEN => wen_a28,
         C_BLK => cblk,
         C_WIDTH => width28,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_28);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_27 : RAM64x18 
      PORT MAP (
         A_DOUT => readData27,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr27,
         B_ADDR => readAddr27,
         A_WIDTH => width27,
         B_WIDTH => width27,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr27,
         C_DIN => writeData27,
         C_WEN => wen_a27,
         C_BLK => cblk,
         C_WIDTH => width27,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_27);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_26 : RAM64x18 
      PORT MAP (
         A_DOUT => readData26,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr26,
         B_ADDR => readAddr26,
         A_WIDTH => width26,
         B_WIDTH => width26,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr26,
         C_DIN => writeData26,
         C_WEN => wen_a26,
         C_BLK => cblk,
         C_WIDTH => width26,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_26);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_25 : RAM64x18 
      PORT MAP (
         A_DOUT => readData25,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr25,
         B_ADDR => readAddr25,
         A_WIDTH => width25,
         B_WIDTH => width25,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr25,
         C_DIN => writeData25,
         C_WEN => wen_a25,
         C_BLK => cblk,
         C_WIDTH => width25,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_25);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_24 : RAM64x18 
      PORT MAP (
         A_DOUT => readData24,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr24,
         B_ADDR => readAddr24,
         A_WIDTH => width24,
         B_WIDTH => width24,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr24,
         C_DIN => writeData24,
         C_WEN => wen_a24,
         C_BLK => cblk,
         C_WIDTH => width24,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_24);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_23 : RAM64x18 
      PORT MAP (
         A_DOUT => readData23,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr23,
         B_ADDR => readAddr23,
         A_WIDTH => width23,
         B_WIDTH => width23,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr23,
         C_DIN => writeData23,
         C_WEN => wen_a23,
         C_BLK => cblk,
         C_WIDTH => width23,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_23);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_22 : RAM64x18 
      PORT MAP (
         A_DOUT => readData22,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr22,
         B_ADDR => readAddr22,
         A_WIDTH => width22,
         B_WIDTH => width22,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr22,
         C_DIN => writeData22,
         C_WEN => wen_a22,
         C_BLK => cblk,
         C_WIDTH => width22,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_22);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_21 : RAM64x18 
      PORT MAP (
         A_DOUT => readData21,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr21,
         B_ADDR => readAddr21,
         A_WIDTH => width21,
         B_WIDTH => width21,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr21,
         C_DIN => writeData21,
         C_WEN => wen_a21,
         C_BLK => cblk,
         C_WIDTH => width21,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_21);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_20 : RAM64x18 
      PORT MAP (
         A_DOUT => readData20,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr20,
         B_ADDR => readAddr20,
         A_WIDTH => width20,
         B_WIDTH => width20,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr20,
         C_DIN => writeData20,
         C_WEN => wen_a20,
         C_BLK => cblk,
         C_WIDTH => width20,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_20);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_19 : RAM64x18 
      PORT MAP (
         A_DOUT => readData19,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr19,
         B_ADDR => readAddr19,
         A_WIDTH => width19,
         B_WIDTH => width19,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr19,
         C_DIN => writeData19,
         C_WEN => wen_a19,
         C_BLK => cblk,
         C_WIDTH => width19,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_19);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_18 : RAM64x18 
      PORT MAP (
         A_DOUT => readData18,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr18,
         B_ADDR => readAddr18,
         A_WIDTH => width18,
         B_WIDTH => width18,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr18,
         C_DIN => writeData18,
         C_WEN => wen_a18,
         C_BLK => cblk,
         C_WIDTH => width18,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_18);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_17 : RAM64x18 
      PORT MAP (
         A_DOUT => readData17,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr17,
         B_ADDR => readAddr17,
         A_WIDTH => width17,
         B_WIDTH => width17,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr17,
         C_DIN => writeData17,
         C_WEN => wen_a17,
         C_BLK => cblk,
         C_WIDTH => width17,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_17);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_16 : RAM64x18 
      PORT MAP (
         A_DOUT => readData16,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr16,
         B_ADDR => readAddr16,
         A_WIDTH => width16,
         B_WIDTH => width16,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr16,
         C_DIN => writeData16,
         C_WEN => wen_a16,
         C_BLK => cblk,
         C_WIDTH => width16,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_16);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_15 : RAM64x18 
      PORT MAP (
         A_DOUT => readData15,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr15,
         B_ADDR => readAddr15,
         A_WIDTH => width15,
         B_WIDTH => width15,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr15,
         C_DIN => writeData15,
         C_WEN => wen_a15,
         C_BLK => cblk,
         C_WIDTH => width15,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_15);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_14 : RAM64x18 
      PORT MAP (
         A_DOUT => readData14,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr14,
         B_ADDR => readAddr14,
         A_WIDTH => width14,
         B_WIDTH => width14,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr14,
         C_DIN => writeData14,
         C_WEN => wen_a14,
         C_BLK => cblk,
         C_WIDTH => width14,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_14);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_13 : RAM64x18 
      PORT MAP (
         A_DOUT => readData13,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr13,
         B_ADDR => readAddr13,
         A_WIDTH => width13,
         B_WIDTH => width13,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr13,
         C_DIN => writeData13,
         C_WEN => wen_a13,
         C_BLK => cblk,
         C_WIDTH => width13,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_13);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_12 : RAM64x18 
      PORT MAP (
         A_DOUT => readData12,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr12,
         B_ADDR => readAddr12,
         A_WIDTH => width12,
         B_WIDTH => width12,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr12,
         C_DIN => writeData12,
         C_WEN => wen_a12,
         C_BLK => cblk,
         C_WIDTH => width12,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_12);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_11 : RAM64x18 
      PORT MAP (
         A_DOUT => readData11,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr11,
         B_ADDR => readAddr11,
         A_WIDTH => width11,
         B_WIDTH => width11,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr11,
         C_DIN => writeData11,
         C_WEN => wen_a11,
         C_BLK => cblk,
         C_WIDTH => width11,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_11);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_10 : RAM64x18 
      PORT MAP (
         A_DOUT => readData10,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr10,
         B_ADDR => readAddr10,
         A_WIDTH => width10,
         B_WIDTH => width10,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr10,
         C_DIN => writeData10,
         C_WEN => wen_a10,
         C_BLK => cblk,
         C_WIDTH => width10,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_10);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_9 : RAM64x18 
      PORT MAP (
         A_DOUT => readData9,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr9,
         B_ADDR => readAddr9,
         A_WIDTH => width9,
         B_WIDTH => width9,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr9,
         C_DIN => writeData9,
         C_WEN => wen_a9,
         C_BLK => cblk,
         C_WIDTH => width9,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_9);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_8 : RAM64x18 
      PORT MAP (
         A_DOUT => readData8,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr8,
         B_ADDR => readAddr8,
         A_WIDTH => width8,
         B_WIDTH => width8,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr8,
         C_DIN => writeData8,
         C_WEN => wen_a8,
         C_BLK => cblk,
         C_WIDTH => width8,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_8);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_7 : RAM64x18 
      PORT MAP (
         A_DOUT => readData7,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr7,
         B_ADDR => readAddr7,
         A_WIDTH => width7,
         B_WIDTH => width7,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr7,
         C_DIN => writeData7,
         C_WEN => wen_a7,
         C_BLK => cblk,
         C_WIDTH => width7,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_7);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_6 : RAM64x18 
      PORT MAP (
         A_DOUT => readData6,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr6,
         B_ADDR => readAddr6,
         A_WIDTH => width6,
         B_WIDTH => width6,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr6,
         C_DIN => writeData6,
         C_WEN => wen_a6,
         C_BLK => cblk,
         C_WIDTH => width6,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_6);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_5 : RAM64x18 
      PORT MAP (
         A_DOUT => readData5,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr5,
         B_ADDR => readAddr5,
         A_WIDTH => width5,
         B_WIDTH => width5,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr5,
         C_DIN => writeData5,
         C_WEN => wen_a5,
         C_BLK => cblk,
         C_WIDTH => width5,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_5);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_4 : RAM64x18 
      PORT MAP (
         A_DOUT => readData4,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr4,
         B_ADDR => readAddr4,
         A_WIDTH => width4,
         B_WIDTH => width4,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr4,
         C_DIN => writeData4,
         C_WEN => wen_a4,
         C_BLK => cblk,
         C_WIDTH => width4,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_4);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_3 : RAM64x18 
      PORT MAP (
         A_DOUT => readData3,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr3,
         B_ADDR => readAddr3,
         A_WIDTH => width3,
         B_WIDTH => width3,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr3,
         C_DIN => writeData3,
         C_WEN => wen_a3,
         C_BLK => cblk,
         C_WIDTH => width3,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_3);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_2 : RAM64x18 
      PORT MAP (
         A_DOUT => readData2,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr2,
         B_ADDR => readAddr2,
         A_WIDTH => width2,
         B_WIDTH => width2,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr2,
         C_DIN => writeData2,
         C_WEN => wen_a2,
         C_BLK => cblk,
         C_WIDTH => width2,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_2);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_1 : RAM64x18 
      PORT MAP (
         A_DOUT => readData1,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr1,
         B_ADDR => readAddr1,
         A_WIDTH => width1,
         B_WIDTH => width1,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr1,
         C_DIN => writeData1,
         C_WEN => wen_a1,
         C_BLK => cblk,
         C_WIDTH => width1,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_1);   
   
   
   --                    .A_BLK(2'b11),                 .B_BLK(2'b11),
   block_0 : RAM64x18 
      PORT MAP (
         A_DOUT => readData0,
         B_DOUT => open,
         A_ADDR_CLK => '1',
         B_ADDR_CLK => '1',
         A_ADDR_EN => '1',
         B_ADDR_EN => '1',
         A_ADDR_LAT => '1',
         B_ADDR_LAT => '1',
         A_ADDR_ARST_N => resetn,
         B_ADDR_ARST_N => resetn,
         A_ADDR_SRST_N => '1',
         B_ADDR_SRST_N => '1',
         A_DOUT_CLK => clk,
         B_DOUT_CLK => clk,
         A_DOUT_EN => '1',
         B_DOUT_EN => '1',
         A_DOUT_LAT => '0',
         B_DOUT_LAT => '0',
         A_DOUT_ARST_N => resetn,
         B_DOUT_ARST_N => resetn,
         A_DOUT_SRST_N => '1',
         B_DOUT_SRST_N => '1',
         A_ADDR => readAddr0,
         B_ADDR => readAddr0,
         A_WIDTH => width0,
         B_WIDTH => width0,
         A_BLK => ablk,
         B_BLK => bblk,
         A_EN => '1',
         B_EN => '1',
         C_CLK => clk,
         C_ADDR => writeAddr0,
         C_DIN => writeData0,
         C_WEN => wen_a0,
         C_BLK => cblk,
         C_WIDTH => width0,
         C_EN => '1',
         SII_LOCK => '0',
         BUSY => u_BUSY_0);   
   
   u_4K_BUSY_all_xhdl2 <= u_BUSY_0 OR u_BUSY_1 OR u_BUSY_2 OR u_BUSY_3 OR 
   u_BUSY_4 OR u_BUSY_5 OR u_BUSY_6 OR u_BUSY_7 OR u_BUSY_8 OR u_BUSY_9 
   OR u_BUSY_10 OR u_BUSY_11 OR u_BUSY_12 OR u_BUSY_13 OR u_BUSY_14 OR 
   u_BUSY_15 OR u_BUSY_16 OR u_BUSY_17 OR u_BUSY_18 OR u_BUSY_19 OR 
   u_BUSY_20 OR u_BUSY_21 OR u_BUSY_22 OR u_BUSY_23 OR u_BUSY_24 OR 
   u_BUSY_25 OR u_BUSY_26 OR u_BUSY_27 OR u_BUSY_28 OR u_BUSY_29 OR 
   u_BUSY_30 OR u_BUSY_31 OR u_BUSY_32 OR u_BUSY_33 OR u_BUSY_34 OR 
   u_BUSY_35 OR u_BUSY_36 OR u_BUSY_37 OR u_BUSY_38 OR u_BUSY_39 OR 
   u_BUSY_40 OR u_BUSY_41 OR u_BUSY_42 OR u_BUSY_43 OR u_BUSY_44 OR 
   u_BUSY_45 OR u_BUSY_46 OR u_BUSY_47 OR u_BUSY_48 OR u_BUSY_49 OR 
   u_BUSY_50 OR u_BUSY_51 OR u_BUSY_52 OR u_BUSY_53 OR u_BUSY_54 OR 
   u_BUSY_55 OR u_BUSY_56 OR u_BUSY_57 OR u_BUSY_58 OR u_BUSY_59 OR 
   u_BUSY_60 OR u_BUSY_61 OR u_BUSY_62 OR u_BUSY_63 OR u_BUSY_64 OR 
   u_BUSY_65 OR u_BUSY_66 OR u_BUSY_67 OR u_BUSY_68 OR u_BUSY_69 OR 
   u_BUSY_70 OR u_BUSY_71 ;

END ARCHITECTURE translated;
