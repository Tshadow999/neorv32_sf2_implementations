----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Fri Oct 18 08:59:04 2024
-- Parameters for COREAXI
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant ADDR_HGS_CFG : integer := 1;
    constant AXI_DWIDTH : integer := 64;
    constant FAMILY : integer := 24;
    constant FEED_THROUGH : 
    constant HDL_License : string( 1 to 1 ) := "U";
    constant HGS_CFG : integer := 1;
    constant ID_WIDTH : integer := 4;
    constant INP_REG_BUF : integer := 1;
    constant M0_SLAVE0ENABLE : integer := 1;
    constant M0_SLAVE1ENABLE : integer := 0;
    constant M0_SLAVE2ENABLE : integer := 0;
    constant M0_SLAVE3ENABLE : integer := 0;
    constant M0_SLAVE4ENABLE : integer := 0;
    constant M0_SLAVE5ENABLE : integer := 0;
    constant M0_SLAVE6ENABLE : integer := 0;
    constant M0_SLAVE7ENABLE : integer := 0;
    constant M0_SLAVE8ENABLE : integer := 0;
    constant M0_SLAVE9ENABLE : integer := 0;
    constant M0_SLAVE10ENABLE : integer := 0;
    constant M0_SLAVE11ENABLE : integer := 0;
    constant M0_SLAVE12ENABLE : integer := 0;
    constant M0_SLAVE13ENABLE : integer := 0;
    constant M0_SLAVE14ENABLE : integer := 0;
    constant M0_SLAVE15ENABLE : integer := 0;
    constant M0_SLAVE16ENABLE : integer := 0;
    constant M1_SLAVE0ENABLE : integer := 0;
    constant M1_SLAVE1ENABLE : integer := 0;
    constant M1_SLAVE2ENABLE : integer := 0;
    constant M1_SLAVE3ENABLE : integer := 0;
    constant M1_SLAVE4ENABLE : integer := 0;
    constant M1_SLAVE5ENABLE : integer := 0;
    constant M1_SLAVE6ENABLE : integer := 0;
    constant M1_SLAVE7ENABLE : integer := 0;
    constant M1_SLAVE8ENABLE : integer := 0;
    constant M1_SLAVE9ENABLE : integer := 0;
    constant M1_SLAVE10ENABLE : integer := 0;
    constant M1_SLAVE11ENABLE : integer := 0;
    constant M1_SLAVE12ENABLE : integer := 0;
    constant M1_SLAVE13ENABLE : integer := 0;
    constant M1_SLAVE14ENABLE : integer := 0;
    constant M1_SLAVE15ENABLE : integer := 0;
    constant M1_SLAVE16ENABLE : integer := 0;
    constant M2_SLAVE0ENABLE : integer := 0;
    constant M2_SLAVE1ENABLE : integer := 0;
    constant M2_SLAVE2ENABLE : integer := 0;
    constant M2_SLAVE3ENABLE : integer := 0;
    constant M2_SLAVE4ENABLE : integer := 0;
    constant M2_SLAVE5ENABLE : integer := 0;
    constant M2_SLAVE6ENABLE : integer := 0;
    constant M2_SLAVE7ENABLE : integer := 0;
    constant M2_SLAVE8ENABLE : integer := 0;
    constant M2_SLAVE9ENABLE : integer := 0;
    constant M2_SLAVE10ENABLE : integer := 0;
    constant M2_SLAVE11ENABLE : integer := 0;
    constant M2_SLAVE12ENABLE : integer := 0;
    constant M2_SLAVE13ENABLE : integer := 0;
    constant M2_SLAVE14ENABLE : integer := 0;
    constant M2_SLAVE15ENABLE : integer := 0;
    constant M2_SLAVE16ENABLE : integer := 0;
    constant M3_SLAVE0ENABLE : integer := 0;
    constant M3_SLAVE1ENABLE : integer := 0;
    constant M3_SLAVE2ENABLE : integer := 0;
    constant M3_SLAVE3ENABLE : integer := 0;
    constant M3_SLAVE4ENABLE : integer := 0;
    constant M3_SLAVE5ENABLE : integer := 0;
    constant M3_SLAVE6ENABLE : integer := 0;
    constant M3_SLAVE7ENABLE : integer := 0;
    constant M3_SLAVE8ENABLE : integer := 0;
    constant M3_SLAVE9ENABLE : integer := 0;
    constant M3_SLAVE10ENABLE : integer := 0;
    constant M3_SLAVE11ENABLE : integer := 0;
    constant M3_SLAVE12ENABLE : integer := 0;
    constant M3_SLAVE13ENABLE : integer := 0;
    constant M3_SLAVE14ENABLE : integer := 0;
    constant M3_SLAVE15ENABLE : integer := 0;
    constant M3_SLAVE16ENABLE : integer := 0;
    constant MEMSPACE : integer := 3;
    constant NUM_MASTER_SLOT : integer := 1;
    constant OUT_REG_BUF : integer := 1;
    constant RD_ACCEPTANCE : integer := 4;
    constant SC_0 : integer := 0;
    constant SC_1 : integer := 0;
    constant SC_2 : integer := 0;
    constant SC_3 : integer := 0;
    constant SC_4 : integer := 0;
    constant SC_5 : integer := 0;
    constant SC_6 : integer := 0;
    constant SC_7 : integer := 0;
    constant SC_8 : integer := 0;
    constant SC_9 : integer := 0;
    constant SC_10 : integer := 0;
    constant SC_11 : integer := 0;
    constant SC_12 : integer := 0;
    constant SC_13 : integer := 0;
    constant SC_14 : integer := 0;
    constant SC_15 : integer := 0;
    constant testbench : string( 1 to 4 ) := "USER";
end coreparameters;
